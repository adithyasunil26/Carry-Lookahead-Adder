* SPICE3 file created from nor.ext - technology: scmos
.include ../TSMC_180nm.txt
* D G S B
.param SUPPLY=1.8V
.param LAMBDA=0.09u
.param length={2*LAMBDA}
.param w={6*LAMBDA}
.global gnd vdd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

va a gnd pulse 1.8 0 0ns 10ps 10ps 10ns 20ns
vb b gnd pulse 1.8 0 0ns 10ps 10ps 20ns 40ns

M1000 out b a_13_6# w_0_0# CMOSP w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1001 a_13_6# a vdd w_0_0# CMOSP w=24 l=2
+  ad=0 pd=0 as=120 ps=58
M1002 gnd b out Gnd CMOSN w=6 l=2
+  ad=60 pd=44 as=48 ps=28
M1003 out a gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out w_0_0# 0.05fF
C1 b a 0.24fF
C2 gnd a 0.05fF
C3 vdd w_0_0# 0.08fF
C4 b w_0_0# 0.06fF
C5 a w_0_0# 0.06fF
C6 out vdd 0.03fF
C7 out b 0.16fF
C8 gnd out 0.18fF
C9 out a 0.02fF
C10 gnd Gnd 0.13fF
C11 out Gnd 0.09fF
C12 vdd Gnd 0.05fF
C13 b Gnd 0.20fF
C14 a Gnd 0.18fF
C15 w_0_0# Gnd 1.23fF

.tran 100p 40n

.control
set hcopypscolor = 0
set color0=white 
set color1=black 

run
set curplottitle="Adithya-2019102005-nand-layout"

hardcopy nor.eps v(a)+4 v(b)+2 v(out)
.endc
