* SPICE3 file created from ckt.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 gnd ffi_0/q inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in ffi_0/q nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd ffi_0/q inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in ffi_0/q nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1067 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1068 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a gnd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1071 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1072 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op gnd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1074 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1075 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1076 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1078 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1079 gnd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1080 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a gnd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1083 gnd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1084 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b gnd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1086 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1087 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1088 sumffo_0/ffo_0/nand_7/a clk gnd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1090 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1091 gnd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1092 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a gnd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1095 gnd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1096 z1o sumffo_0/ffo_0/nand_7/a gnd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1098 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1099 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1101 sumffo_0/ffo_0/nand_0/b clk gnd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1102 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_0/xor_0/inv_1/op ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_0/xor_0/inv_1/op ffi_0/q gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 gnd ffi_0/q sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 sumffo_0/ffo_0/d ffi_0/q sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1115 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1116 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a gnd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1119 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1120 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op gnd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1122 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1123 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1124 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1127 gnd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1128 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a gnd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1130 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1131 gnd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1132 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b gnd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1134 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1135 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1136 sumffo_2/ffo_0/nand_7/a clk gnd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1139 gnd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1140 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a gnd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1143 gnd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1144 z3o sumffo_2/ffo_0/nand_7/a gnd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1146 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1147 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 sumffo_2/ffo_0/nand_0/b clk gnd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1153 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1154 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1155 sumffo_2/ffo_0/d ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1156 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1157 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1158 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1163 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1164 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a gnd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1166 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1167 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1168 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op gnd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1170 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1171 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1172 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a gnd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1179 gnd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1180 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b gnd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1183 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1184 sumffo_1/ffo_0/nand_7/a clk gnd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1186 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1187 gnd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1188 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a gnd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1190 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1191 gnd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1192 z2o sumffo_1/ffo_0/nand_7/a gnd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1194 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1195 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 sumffo_1/ffo_0/nand_0/b clk gnd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1211 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1212 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a gnd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1214 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op gnd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1219 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1220 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1223 gnd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1224 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a gnd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1226 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1227 gnd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1228 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b gnd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1230 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1231 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1232 sumffo_3/ffo_0/nand_7/a clk gnd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1235 gnd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1236 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a gnd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1238 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1239 gnd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1240 z4o sumffo_3/ffo_0/nand_7/a gnd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1245 sumffo_3/ffo_0/nand_0/b clk gnd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1246 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1247 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1248 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1249 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1250 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1251 sumffo_3/ffo_0/d ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1252 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1253 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1254 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1259 gnd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1260 ffo_0/nand_3/b ffo_0/nand_1/a gnd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1262 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1263 gnd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1264 ffo_0/nand_1/a ffo_0/inv_0/op gnd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1266 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1267 gnd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1268 ffo_0/nand_3/a ffo_0/d gnd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1270 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1271 gnd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1272 ffo_0/nand_1/b ffo_0/nand_3/a gnd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1274 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1275 gnd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1276 ffo_0/nand_6/a ffo_0/nand_3/b gnd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1278 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1279 gnd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1280 ffo_0/nand_7/a clk gnd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1282 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1283 gnd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1284 ffo_0/qbar ffo_0/nand_6/a gnd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1286 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1287 gnd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1288 couto ffo_0/nand_7/a gnd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffo_0/inv_0/op ffo_0/d gnd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1293 ffo_0/nand_0/b clk gnd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1294 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1295 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1297 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1298 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1299 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1301 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1303 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1305 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1306 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1307 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1309 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1311 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1313 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1314 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1315 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1317 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1318 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1319 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1320 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1321 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1323 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1325 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1327 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1329 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1330 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1331 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipg_0/pggen_0/nand_0/a_13_n26# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 gnd ffipg_0/ffi_0/q cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 cla_0/g0 ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 cla_0/g0 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1337 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1338 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1339 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 gnd ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1341 ffipg_0/k ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1342 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1343 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1344 ffipg_0/pggen_0/xor_0/a_10_n43# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 nor_0/a ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1349 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 gnd ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1351 nor_0/a ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 ffipg_0/ffi_0/nand_1/a_13_n26# ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/a gnd ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipg_0/ffi_0/nand_0/a_13_n26# ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 gnd clk ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/inv_0/op gnd ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 ffipg_0/ffi_0/nand_1/a clk ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1361 gnd clk ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1362 ffipg_0/ffi_0/nand_3/a y1in gnd ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 ffipg_0/ffi_0/nand_3/a clk ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipg_0/ffi_0/nand_3/a_13_n26# ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 gnd ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/a gnd ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipg_0/ffi_0/nand_4/a_13_n26# ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1369 gnd ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1370 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_3/b gnd ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1371 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 ffipg_0/ffi_0/nand_5/a_13_n26# ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1373 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1374 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/inv_1/op gnd ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1376 ffipg_0/ffi_0/nand_6/a_13_n26# ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1377 gnd ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1378 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/a gnd ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1380 ffipg_0/ffi_0/nand_7/a_13_n26# ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1381 gnd ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1382 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a gnd ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1384 ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1385 ffipg_0/ffi_0/inv_0/op y1in gnd ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1386 ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1387 ffipg_0/ffi_0/inv_1/op clk gnd ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipg_0/ffi_1/nand_1/a_13_n26# ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a gnd ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipg_0/ffi_1/nand_0/a_13_n26# ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 gnd clk ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/inv_0/op gnd ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipg_0/ffi_1/nand_1/a clk ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 gnd clk ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipg_0/ffi_1/nand_3/a x1in gnd ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipg_0/ffi_1/nand_3/a clk ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipg_0/ffi_1/nand_3/a_13_n26# ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 gnd ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/a gnd ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipg_0/ffi_1/nand_4/a_13_n26# ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 gnd ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_3/b gnd ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipg_0/ffi_1/nand_5/a_13_n26# ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/inv_1/op gnd ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipg_0/ffi_1/nand_6/a_13_n26# ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 gnd ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/a gnd ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipg_0/ffi_1/nand_7/a_13_n26# ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1417 gnd ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1418 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a gnd ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1421 ffipg_0/ffi_1/inv_0/op x1in gnd ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1422 ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1423 ffipg_0/ffi_1/inv_1/op clk gnd ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1425 ffo_0/d inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1426 ffipg_1/pggen_0/nand_0/a_13_n26# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1427 gnd ffipg_1/ffi_0/q cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 cla_0/l ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 cla_0/l ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1431 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1433 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1434 gnd ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1435 ffipg_1/k ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1436 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1437 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1438 ffipg_1/pggen_0/xor_0/a_10_n43# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 cla_1/p0 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1443 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 gnd ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1445 cla_1/p0 ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 ffipg_1/ffi_0/nand_1/a_13_n26# ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1447 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1448 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a gnd ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1450 ffipg_1/ffi_0/nand_0/a_13_n26# ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1451 gnd clk ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1452 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/inv_0/op gnd ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 ffipg_1/ffi_0/nand_1/a clk ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1455 gnd clk ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1456 ffipg_1/ffi_0/nand_3/a y2in gnd ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 ffipg_1/ffi_0/nand_3/a clk ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1458 ffipg_1/ffi_0/nand_3/a_13_n26# ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1459 gnd ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1460 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/a gnd ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 ffipg_1/ffi_0/nand_4/a_13_n26# ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1463 gnd ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1464 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_3/b gnd ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1466 ffipg_1/ffi_0/nand_5/a_13_n26# ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1467 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1468 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/inv_1/op gnd ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1470 ffipg_1/ffi_0/nand_6/a_13_n26# ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 gnd ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a gnd ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 ffipg_1/ffi_0/nand_7/a_13_n26# ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 gnd ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a gnd ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 ffipg_1/ffi_0/inv_0/op y2in gnd ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1480 ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1481 ffipg_1/ffi_0/inv_1/op clk gnd ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 ffipg_1/ffi_1/nand_1/a_13_n26# ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a gnd ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 ffipg_1/ffi_1/nand_0/a_13_n26# ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 gnd clk ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/inv_0/op gnd ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 ffipg_1/ffi_1/nand_1/a clk ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 gnd clk ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 ffipg_1/ffi_1/nand_3/a x2in gnd ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 ffipg_1/ffi_1/nand_3/a clk ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 ffipg_1/ffi_1/nand_3/a_13_n26# ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 gnd ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/a gnd ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 ffipg_1/ffi_1/nand_4/a_13_n26# ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 gnd ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_3/b gnd ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 ffipg_1/ffi_1/nand_5/a_13_n26# ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1503 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1504 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/inv_1/op gnd ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1505 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 ffipg_1/ffi_1/nand_6/a_13_n26# ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1507 gnd ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1508 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a gnd ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 ffipg_1/ffi_1/nand_7/a_13_n26# ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1511 gnd ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1512 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a gnd ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1513 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1514 ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1515 ffipg_1/ffi_1/inv_0/op x2in gnd ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1516 ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1517 ffipg_1/ffi_1/inv_1/op clk gnd ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1518 ffipg_2/pggen_0/nand_0/a_13_n26# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 gnd ffipg_2/ffi_0/q cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1520 cla_0/l ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 cla_0/l ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1523 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1524 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1525 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 gnd ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1527 ffipg_2/k ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1528 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1529 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1530 ffipg_2/pggen_0/xor_0/a_10_n43# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1534 cla_2/p0 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1535 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 gnd ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1537 cla_2/p0 ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 ffipg_2/ffi_0/nand_1/a_13_n26# ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a gnd ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 ffipg_2/ffi_0/nand_0/a_13_n26# ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 gnd clk ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/inv_0/op gnd ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 ffipg_2/ffi_0/nand_1/a clk ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 gnd clk ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 ffipg_2/ffi_0/nand_3/a y3in gnd ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 ffipg_2/ffi_0/nand_3/a clk ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 ffipg_2/ffi_0/nand_3/a_13_n26# ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1551 gnd ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1552 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/a gnd ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 ffipg_2/ffi_0/nand_4/a_13_n26# ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1555 gnd ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1556 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_3/b gnd ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 ffipg_2/ffi_0/nand_5/a_13_n26# ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1559 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1560 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/inv_1/op gnd ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1561 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1562 ffipg_2/ffi_0/nand_6/a_13_n26# ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1563 gnd ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1564 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/a gnd ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1566 ffipg_2/ffi_0/nand_7/a_13_n26# ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 gnd ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a gnd ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1571 ffipg_2/ffi_0/inv_0/op y3in gnd ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1572 ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1573 ffipg_2/ffi_0/inv_1/op clk gnd ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 ffipg_2/ffi_1/nand_1/a_13_n26# ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a gnd ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 ffipg_2/ffi_1/nand_0/a_13_n26# ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 gnd clk ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/inv_0/op gnd ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 ffipg_2/ffi_1/nand_1/a clk ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 gnd clk ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 ffipg_2/ffi_1/nand_3/a x3in gnd ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 ffipg_2/ffi_1/nand_3/a clk ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 ffipg_2/ffi_1/nand_3/a_13_n26# ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 gnd ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/a gnd ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 ffipg_2/ffi_1/nand_4/a_13_n26# ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 gnd ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_3/b gnd ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 ffipg_2/ffi_1/nand_5/a_13_n26# ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/inv_1/op gnd ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 ffipg_2/ffi_1/nand_6/a_13_n26# ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1599 gnd ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1600 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/a gnd ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1601 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 ffipg_2/ffi_1/nand_7/a_13_n26# ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1603 gnd ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1604 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a gnd ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1605 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1607 ffipg_2/ffi_1/inv_0/op x3in gnd ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1608 ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1609 ffipg_2/ffi_1/inv_1/op clk gnd ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1610 ffi_0/nand_1/a_13_n26# ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1611 gnd ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1612 ffi_0/nand_3/b ffi_0/nand_1/a gnd ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1614 ffi_0/nand_0/a_13_n26# ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 gnd clk ffi_0/nand_1/a ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 ffi_0/nand_1/a ffi_0/inv_0/op gnd ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 ffi_0/nand_1/a clk ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 gnd clk ffi_0/nand_3/a ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 ffi_0/nand_3/a cinin gnd ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 ffi_0/nand_3/a clk ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 ffi_0/nand_3/a_13_n26# ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 gnd ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 ffi_0/nand_1/b ffi_0/nand_3/a gnd ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 ffi_0/nand_4/a_13_n26# ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 gnd ffi_0/inv_1/op ffi_0/nand_6/a ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 ffi_0/nand_6/a ffi_0/nand_3/b gnd ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 ffi_0/nand_6/a ffi_0/inv_1/op ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 ffi_0/nand_5/a_13_n26# ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 gnd ffi_0/nand_1/b ffi_0/nand_7/a ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 ffi_0/nand_7/a ffi_0/inv_1/op gnd ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 ffi_0/nand_7/a ffi_0/nand_1/b ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 ffi_0/nand_6/a_13_n26# ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 gnd ffi_0/q nor_0/b ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 nor_0/b ffi_0/nand_6/a gnd ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 nor_0/b ffi_0/q ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 ffi_0/nand_7/a_13_n26# ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 gnd nor_0/b ffi_0/q ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 ffi_0/q ffi_0/nand_7/a gnd ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 ffi_0/q nor_0/b ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1643 ffi_0/inv_0/op cinin gnd ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1644 ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1645 ffi_0/inv_1/op clk gnd ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 ffipg_3/pggen_0/nand_0/a_13_n26# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1647 gnd ffipg_3/ffi_0/q cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1648 cla_2/g1 ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1649 cla_2/g1 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 gnd ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 ffipg_3/k ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 ffipg_3/pggen_0/xor_0/a_10_n43# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 cla_2/p1 ffipg_3/ffi_1/q ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1663 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 gnd ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1665 cla_2/p1 ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1666 ffipg_3/ffi_0/nand_1/a_13_n26# ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/a gnd ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffipg_3/ffi_0/nand_0/a_13_n26# ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 gnd clk ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/inv_0/op gnd ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffipg_3/ffi_0/nand_1/a clk ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 gnd clk ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffipg_3/ffi_0/nand_3/a y4in gnd ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffipg_3/ffi_0/nand_3/a clk ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffipg_3/ffi_0/nand_3/a_13_n26# ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 gnd ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/a gnd ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffipg_3/ffi_0/nand_4/a_13_n26# ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 gnd ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_3/b gnd ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffipg_3/ffi_0/nand_5/a_13_n26# ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/inv_1/op gnd ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffipg_3/ffi_0/nand_6/a_13_n26# ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 gnd ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/a gnd ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffipg_3/ffi_0/nand_7/a_13_n26# ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1695 gnd ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1696 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a gnd ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1697 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 ffipg_3/ffi_0/inv_0/op y4in gnd ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 ffipg_3/ffi_0/inv_1/op clk gnd ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 ffipg_3/ffi_1/nand_1/a_13_n26# ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1703 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1704 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/a gnd ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1705 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1706 ffipg_3/ffi_1/nand_0/a_13_n26# ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1707 gnd clk ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1708 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/inv_0/op gnd ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1709 ffipg_3/ffi_1/nand_1/a clk ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1711 gnd clk ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1712 ffipg_3/ffi_1/nand_3/a x4in gnd ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1713 ffipg_3/ffi_1/nand_3/a clk ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1714 ffipg_3/ffi_1/nand_3/a_13_n26# ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1715 gnd ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1716 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/a gnd ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1717 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1718 ffipg_3/ffi_1/nand_4/a_13_n26# ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1719 gnd ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1720 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_3/b gnd ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1721 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 ffipg_3/ffi_1/nand_5/a_13_n26# ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1723 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1724 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/inv_1/op gnd ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1725 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1726 ffipg_3/ffi_1/nand_6/a_13_n26# ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1727 gnd ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1728 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/a gnd ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1730 ffipg_3/ffi_1/nand_7/a_13_n26# ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1731 gnd ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1732 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a gnd ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 ffipg_3/ffi_1/inv_0/op x4in gnd ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffipg_3/ffi_1/inv_1/op clk gnd ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 clk ffo_0/nand_1/b 0.45fF
C1 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C2 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/q 0.31fF
C3 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C4 sumffo_3/ffo_0/nand_6/a gnd 0.33fF
C5 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C6 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C7 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C8 ffipg_2/k nand_2/b 0.06fF
C9 ffipg_3/ffi_0/inv_0/op ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C10 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C11 inv_1/in cla_0/n 0.02fF
C12 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C13 cla_0/inv_0/op gnd 0.27fF
C14 ffi_0/nand_6/w_0_0# gnd 0.10fF
C15 cla_0/g0 ffipg_1/k 0.06fF
C16 ffi_0/nand_1/a ffi_0/nand_1/w_0_0# 0.06fF
C17 ffipg_2/ffi_1/nand_7/w_0_0# ffipg_2/ffi_1/nand_7/a 0.06fF
C18 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_3/b 0.04fF
C19 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a 0.31fF
C20 nor_0/b ffi_0/nand_6/a 0.00fF
C21 ffo_0/nand_6/a ffo_0/nand_6/w_0_0# 0.06fF
C22 clk sumffo_2/ffo_0/d 0.25fF
C23 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op 0.13fF
C24 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d 0.04fF
C25 gnd ffipg_0/ffi_1/nand_6/w_0_0# 0.10fF
C26 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C27 gnd inv_8/in 0.43fF
C28 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/a 0.00fF
C29 ffi_0/nand_1/b ffi_0/nand_1/a 0.31fF
C30 clk ffipg_1/ffi_1/nand_3/a 0.13fF
C31 ffipg_1/ffi_0/inv_0/op clk 0.32fF
C32 x3in ffipg_2/ffi_1/inv_1/op 0.01fF
C33 inv_8/w_0_6# inv_8/in 0.10fF
C34 sumffo_1/ffo_0/d gnd 0.41fF
C35 sumffo_2/ffo_0/nand_1/a gnd 0.33fF
C36 cla_0/g0 gnd 1.11fF
C37 cla_2/g1 ffipg_3/ffi_0/q 0.13fF
C38 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C39 sumffo_1/xor_0/inv_0/op ffi_0/q 0.06fF
C40 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C41 nor_0/b ffipg_0/k 0.06fF
C42 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C43 ffipg_1/ffi_1/q ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C44 gnd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C45 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C46 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/k 0.45fF
C47 nor_3/w_0_0# inv_6/in 0.11fF
C48 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C49 clk ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C50 ffipg_2/ffi_1/nand_5/w_0_0# gnd 0.10fF
C51 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# 0.04fF
C52 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b 0.32fF
C53 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/a 0.06fF
C54 ffipg_2/ffi_0/inv_0/op ffipg_2/ffi_0/inv_0/w_0_6# 0.03fF
C55 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C56 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C57 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q 0.27fF
C58 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/b 0.31fF
C59 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_0/inv_1/op 0.75fF
C60 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a 0.31fF
C61 cla_0/g0 inv_0/op 0.33fF
C62 ffipg_3/ffi_1/inv_1/w_0_6# gnd 0.06fF
C63 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C64 gnd ffipg_2/ffi_1/nand_2/w_0_0# 0.10fF
C65 sumffo_3/sbar sumffo_3/ffo_0/nand_7/a 0.31fF
C66 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/ffi_0/q 0.06fF
C67 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/q 0.31fF
C68 ffipg_3/ffi_0/nand_2/w_0_0# ffipg_3/ffi_0/nand_3/a 0.04fF
C69 ffipg_1/pggen_0/xor_0/a_10_10# gnd 0.93fF
C70 ffo_0/qbar ffo_0/nand_6/a 0.00fF
C71 sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d 0.52fF
C72 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/qbar 0.00fF
C73 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/nand_1/b 0.06fF
C74 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/k 0.01fF
C75 cla_0/l cla_1/inv_0/op 0.35fF
C76 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/nand_6/a 0.06fF
C77 y3in ffipg_2/ffi_0/inv_0/op 0.04fF
C78 ffipg_1/ffi_0/nand_3/a clk 0.13fF
C79 ffi_0/nand_6/a gnd 0.33fF
C80 ffipg_0/ffi_0/nand_1/b gnd 0.57fF
C81 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C82 cla_2/p1 cla_2/p0 0.24fF
C83 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/a 0.06fF
C84 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C85 gnd ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C86 ffi_0/nand_3/b ffi_0/nand_1/a 0.00fF
C87 ffipg_1/ffi_1/q ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C88 inv_4/op ffipg_3/k 0.09fF
C89 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_1/b 0.45fF
C90 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C91 gnd ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C92 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C93 gnd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C94 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# 0.04fF
C95 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_3/b 0.04fF
C96 inv_5/in cla_2/l 0.05fF
C97 ffipg_3/ffi_1/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C98 ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C99 sumffo_1/ffo_0/inv_0/w_0_6# gnd 0.06fF
C100 sumffo_0/xor_0/inv_0/op ffi_0/q 0.20fF
C101 nor_2/w_0_0# cla_1/n 0.06fF
C102 ffipg_2/ffi_1/nand_4/w_0_0# ffipg_2/ffi_1/nand_3/b 0.06fF
C103 inv_6/in cla_2/n 0.02fF
C104 ffipg_0/k gnd 0.68fF
C105 ffipg_3/ffi_0/inv_1/op clk 0.07fF
C106 ffipg_2/ffi_1/nand_3/w_0_0# gnd 0.11fF
C107 y1in ffipg_0/ffi_0/inv_1/op 0.01fF
C108 sumffo_3/xor_0/inv_1/op ffi_0/q 0.04fF
C109 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/a 0.06fF
C110 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/inv_0/w_0_6# 0.03fF
C111 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/k 0.02fF
C112 sumffo_3/xor_0/a_10_10# sumffo_3/ffo_0/d 0.45fF
C113 ffi_0/nand_0/a_13_n26# gnd 0.01fF
C114 gnd ffipg_3/ffi_1/nand_3/a 0.33fF
C115 nor_4/b inv_6/in 0.04fF
C116 sumffo_3/xor_0/inv_1/op inv_4/op 0.06fF
C117 ffipg_2/ffi_1/inv_0/op gnd 0.27fF
C118 cla_0/inv_0/op nand_2/b 0.09fF
C119 ffipg_0/ffi_1/q nor_0/a 0.22fF
C120 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C121 ffi_0/nand_0/w_0_0# ffi_0/nand_1/a 0.04fF
C122 ffipg_1/ffi_1/nand_2/w_0_0# x2in 0.06fF
C123 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/a 0.06fF
C124 ffipg_2/ffi_1/q gnd 2.24fF
C125 sumffo_3/ffo_0/nand_5/w_0_0# gnd 0.10fF
C126 y2in clk 0.68fF
C127 ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C128 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C129 clk y4in 0.64fF
C130 cla_2/g1 cla_2/n 0.13fF
C131 ffipg_1/ffi_1/inv_0/w_0_6# x2in 0.06fF
C132 clk sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C133 sumffo_3/ffo_0/nand_3/a gnd 0.33fF
C134 ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# 0.04fF
C135 gnd ffipg_1/ffi_1/qbar 0.67fF
C136 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/d 0.06fF
C137 cla_0/l cla_1/inv_0/in 0.23fF
C138 ffipg_0/ffi_0/inv_0/op y1in 0.04fF
C139 z4o sumffo_3/ffo_0/nand_7/a 0.00fF
C140 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b 0.13fF
C141 cinin ffi_0/inv_0/op 0.04fF
C142 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C143 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_5/w_0_0# 0.04fF
C144 gnd ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C145 sumffo_2/ffo_0/nand_0/w_0_0# gnd 0.10fF
C146 cla_0/g0 nand_2/b 0.13fF
C147 nor_0/b ffi_0/nand_7/a 0.31fF
C148 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C149 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C150 clk ffipg_3/ffi_0/inv_0/op 0.32fF
C151 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C152 gnd ffo_0/inv_1/w_0_6# 0.06fF
C153 cla_1/inv_0/op gnd 0.27fF
C154 ffipg_3/ffi_0/nand_2/w_0_0# gnd 0.10fF
C155 ffipg_2/ffi_1/inv_1/op gnd 1.85fF
C156 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C157 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/qbar 0.31fF
C158 sumffo_0/ffo_0/nand_1/w_0_0# gnd 0.10fF
C159 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a 0.31fF
C160 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C161 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C162 gnd sumffo_2/ffo_0/nand_3/b 0.74fF
C163 clk ffi_0/nand_3/a 0.13fF
C164 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_1/inv_1/op 0.75fF
C165 ffipg_0/ffi_0/nand_0/w_0_0# ffipg_0/ffi_0/nand_1/a 0.04fF
C166 clk sumffo_0/ffo_0/d 0.25fF
C167 ffipg_0/ffi_1/nand_0/w_0_0# ffipg_0/ffi_1/nand_1/a 0.04fF
C168 ffipg_3/ffi_0/nand_4/w_0_0# gnd 0.10fF
C169 nor_3/b inv_6/in 0.16fF
C170 gnd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C171 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C172 sumffo_3/xor_0/a_10_10# gnd 0.93fF
C173 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C174 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C175 sumffo_1/ffo_0/nand_0/b clk 0.04fF
C176 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C177 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/qbar 0.00fF
C178 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/a 0.06fF
C179 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_3/a 0.06fF
C180 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/inv_0/op 0.06fF
C181 gnd ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C182 clk ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C183 ffipg_0/ffi_1/inv_0/op gnd 0.27fF
C184 ffipg_2/ffi_0/nand_2/w_0_0# gnd 0.10fF
C185 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# 0.04fF
C186 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a 0.13fF
C187 sumffo_0/ffo_0/nand_7/w_0_0# z1o 0.04fF
C188 cla_0/nor_1/w_0_0# cla_0/inv_0/in 0.05fF
C189 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_3/b 0.04fF
C190 gnd ffipg_2/ffi_0/nand_1/b 0.57fF
C191 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C192 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/qbar 0.31fF
C193 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/qbar 0.00fF
C194 gnd ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C195 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar 0.32fF
C196 sumffo_0/xor_0/a_10_10# ffi_0/q 0.12fF
C197 x3in gnd 0.22fF
C198 ffipg_0/ffi_1/nand_7/a gnd 0.37fF
C199 ffo_0/nand_1/a gnd 0.33fF
C200 cla_0/nand_0/a_13_n26# gnd 0.00fF
C201 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/w_0_0# 0.04fF
C202 clk ffo_0/nand_4/w_0_0# 0.06fF
C203 ffi_0/nand_1/b ffi_0/inv_1/op 0.45fF
C204 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# 0.04fF
C205 cla_2/p1 cla_2/l 0.02fF
C206 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C207 ffi_0/nand_7/a gnd 0.33fF
C208 sumffo_2/xor_0/w_n3_4# ffi_0/q 0.00fF
C209 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C210 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_0/op 0.06fF
C211 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_1/inv_1/op 0.75fF
C212 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C213 sumffo_0/ffo_0/inv_0/w_0_6# gnd 0.06fF
C214 sumffo_0/ffo_0/nand_1/a gnd 0.44fF
C215 ffi_0/inv_1/op cinin 0.01fF
C216 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C217 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C218 ffo_0/nand_1/b ffo_0/nand_3/b 0.32fF
C219 inv_7/op ffi_0/q 0.31fF
C220 ffi_0/nand_0/w_0_0# ffi_0/inv_0/op 0.06fF
C221 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# 0.04fF
C222 cla_1/inv_0/in gnd 0.34fF
C223 ffipg_2/ffi_0/inv_1/op gnd 1.85fF
C224 ffipg_0/ffi_1/inv_1/op gnd 1.85fF
C225 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C226 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C227 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C228 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/ffi_0/q 0.06fF
C229 cla_1/n nor_2/b 0.39fF
C230 cla_1/nor_0/w_0_0# cla_1/p0 0.06fF
C231 cla_0/l inv_7/in 0.13fF
C232 gnd ffipg_1/ffi_1/nand_0/a_13_n26# 0.01fF
C233 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C234 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C235 ffipg_2/ffi_0/q cla_2/p0 0.03fF
C236 ffipg_1/ffi_1/inv_1/w_0_6# ffipg_1/ffi_1/inv_1/op 0.04fF
C237 gnd ffipg_3/ffi_0/nand_3/a 0.33fF
C238 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_1/b 0.45fF
C239 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C240 ffipg_2/ffi_0/nand_7/w_0_0# gnd 0.10fF
C241 gnd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C242 sumffo_2/ffo_0/nand_2/w_0_0# gnd 0.10fF
C243 gnd cla_2/nor_0/w_0_0# 0.31fF
C244 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C245 cla_0/l gnd 3.05fF
C246 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C247 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C248 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C249 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d 0.04fF
C250 x3in ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C251 ffipg_1/ffi_0/nand_7/w_0_0# ffipg_1/ffi_0/nand_7/a 0.06fF
C252 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b 0.32fF
C253 inv_3/w_0_6# gnd 0.17fF
C254 ffipg_3/ffi_1/nand_2/w_0_0# x4in 0.06fF
C255 nor_0/w_0_0# cla_0/g0 0.06fF
C256 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C257 nor_0/b inv_0/in 0.16fF
C258 ffipg_1/ffi_1/nand_6/a gnd 0.37fF
C259 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/nand_3/b 0.06fF
C260 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C261 clk sumffo_1/ffo_0/nand_6/a 0.13fF
C262 gnd sumffo_2/sbar 0.62fF
C263 sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d 0.06fF
C264 ffipg_3/ffi_1/nand_2/w_0_0# clk 0.06fF
C265 ffi_0/nand_3/b ffi_0/inv_1/op 0.33fF
C266 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C267 nor_0/b gnd 0.74fF
C268 gnd sumffo_3/ffo_0/d 0.41fF
C269 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C270 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_0/q 0.06fF
C271 ffipg_1/ffi_1/nand_4/w_0_0# gnd 0.10fF
C272 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C273 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C274 clk sumffo_1/ffo_0/nand_1/b 0.45fF
C275 nor_1/b inv_2/in 0.04fF
C276 gnd ffipg_1/ffi_0/nand_6/w_0_0# 0.10fF
C277 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C278 gnd ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C279 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C280 nor_4/a gnd 0.40fF
C281 cla_1/l cla_0/l 0.08fF
C282 ffipg_2/k ffipg_2/ffi_0/q 0.07fF
C283 gnd ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C284 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_1/q 0.06fF
C285 inv_8/w_0_6# nor_4/a 0.03fF
C286 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/inv_1/w_0_6# 0.04fF
C287 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a 0.00fF
C288 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/k 0.21fF
C289 gnd sumffo_3/ffo_0/nand_1/w_0_0# 0.10fF
C290 inv_2/in gnd 0.47fF
C291 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C292 cla_1/l inv_3/w_0_6# 0.06fF
C293 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C294 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_1/b 0.04fF
C295 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# 0.04fF
C296 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C297 gnd ffipg_2/ffi_0/nand_5/w_0_0# 0.10fF
C298 clk x1in 0.68fF
C299 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C300 cla_1/inv_0/in cla_1/inv_0/w_0_6# 0.06fF
C301 ffi_0/nand_5/w_0_0# ffi_0/inv_1/op 0.06fF
C302 ffipg_0/ffi_1/qbar gnd 0.67fF
C303 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C304 gnd ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C305 gnd ffipg_1/ffi_0/nand_7/a 0.37fF
C306 sumffo_3/ffo_0/inv_0/op gnd 0.52fF
C307 gnd ffipg_1/k 0.70fF
C308 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C309 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C310 gnd sumffo_0/xor_0/inv_1/op 0.35fF
C311 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C312 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b 0.32fF
C313 ffipg_1/ffi_0/inv_0/op ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C314 nor_4/b inv_9/in 0.16fF
C315 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C316 cla_1/p0 cla_2/p0 0.24fF
C317 gnd inv_0/in 0.30fF
C318 sumffo_3/xor_0/w_n3_4# sumffo_3/ffo_0/d 0.02fF
C319 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/k 0.21fF
C320 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C321 gnd ffipg_3/ffi_0/nand_0/a_13_n26# 0.01fF
C322 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/k 0.01fF
C323 nor_1/b gnd 0.35fF
C324 inv_7/in gnd 0.43fF
C325 gnd ffipg_1/ffi_1/nand_3/b 0.74fF
C326 ffipg_0/ffi_0/nand_7/w_0_0# ffipg_0/ffi_0/nand_7/a 0.06fF
C327 ffipg_1/ffi_1/inv_0/op clk 0.32fF
C328 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C329 clk ffi_0/inv_1/w_0_6# 0.06fF
C330 ffipg_1/ffi_0/inv_1/w_0_6# ffipg_1/ffi_0/inv_1/op 0.04fF
C331 ffo_0/nand_6/a ffo_0/nand_4/w_0_0# 0.04fF
C332 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C333 clk ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C334 gnd sumffo_0/xor_0/inv_1/w_0_6# 0.06fF
C335 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b 0.32fF
C336 sumffo_0/ffo_0/nand_6/a gnd 0.33fF
C337 inv_8/w_0_6# gnd 0.15fF
C338 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C339 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C340 gnd ffipg_3/ffi_1/nand_5/w_0_0# 0.10fF
C341 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/sbar 0.06fF
C342 inv_0/op inv_0/in 0.04fF
C343 gnd ffipg_3/ffi_1/nand_7/a 0.37fF
C344 gnd ffipg_3/ffi_0/nand_7/a 0.37fF
C345 ffipg_1/ffi_0/nand_3/b gnd 0.74fF
C346 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C347 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/q 0.06fF
C348 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a 0.13fF
C349 sumffo_1/xor_0/inv_1/op ffipg_1/k 0.06fF
C350 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C351 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C352 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_1/b 0.45fF
C353 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C354 cla_0/l nand_2/b 0.06fF
C355 nor_4/b nor_4/w_0_0# 0.06fF
C356 sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d 0.06fF
C357 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C358 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# 0.04fF
C359 sumffo_3/ffo_0/nand_0/b clk 0.04fF
C360 ffipg_1/ffi_1/nand_7/a gnd 0.37fF
C361 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/b 0.32fF
C362 inv_0/op gnd 0.27fF
C363 ffipg_1/ffi_1/nand_0/w_0_0# gnd 0.10fF
C364 inv_9/in ffo_0/d 0.04fF
C365 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_7/a 0.04fF
C366 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C367 ffipg_2/k cla_1/p0 0.06fF
C368 inv_3/w_0_6# nand_2/b 0.06fF
C369 gnd ffipg_3/ffi_1/nand_1/a 0.44fF
C370 cla_2/g1 cla_2/inv_0/op 0.35fF
C371 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_3/b 0.33fF
C372 sumffo_1/xor_0/inv_1/op gnd 0.35fF
C373 cla_2/nand_0/w_0_0# gnd 0.18fF
C374 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# 0.04fF
C375 cla_1/l gnd 0.40fF
C376 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/inv_1/op 0.33fF
C377 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a 0.31fF
C378 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/d 0.06fF
C379 sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# 0.04fF
C380 sumffo_3/xor_0/w_n3_4# gnd 0.12fF
C381 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/qbar 0.06fF
C382 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_3/b 0.33fF
C383 ffo_0/nand_7/a gnd 0.33fF
C384 ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.32fF
C385 ffipg_1/ffi_0/q cla_1/p0 0.03fF
C386 ffipg_2/ffi_0/inv_1/w_0_6# clk 0.06fF
C387 gnd ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C388 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C389 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C390 clk x4in 0.68fF
C391 clk ffipg_0/ffi_1/nand_1/a 0.13fF
C392 gnd sumffo_2/xor_0/inv_0/op 0.32fF
C393 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/nand_7/a 0.06fF
C394 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C395 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C396 inv_2/in nand_2/b 0.34fF
C397 ffo_0/d nor_4/w_0_0# 0.03fF
C398 sumffo_0/ffo_0/nand_3/a gnd 0.33fF
C399 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/q 0.04fF
C400 cla_1/inv_0/w_0_6# gnd 0.06fF
C401 ffipg_2/ffi_1/nand_3/a gnd 0.33fF
C402 ffi_0/nand_6/w_0_0# ffi_0/q 0.06fF
C403 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C404 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C405 ffipg_0/ffi_0/q cla_0/g0 0.13fF
C406 clk ffipg_2/ffi_1/nand_1/a 0.13fF
C407 nor_3/b inv_5/w_0_6# 0.17fF
C408 sumffo_3/xor_0/inv_0/op gnd 0.32fF
C409 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/inv_0/w_0_6# 0.03fF
C410 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C411 gnd cla_1/nand_0/w_0_0# 0.10fF
C412 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/b 0.06fF
C413 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C414 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C415 ffi_0/nand_3/w_0_0# ffi_0/nand_3/a 0.06fF
C416 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C417 sumffo_3/ffo_0/nand_7/w_0_0# gnd 0.10fF
C418 inv_8/in ffi_0/q 0.13fF
C419 ffi_0/inv_0/w_0_6# cinin 0.06fF
C420 ffipg_1/k nand_2/b 0.15fF
C421 inv_1/op gnd 0.58fF
C422 ffipg_0/ffi_1/nand_1/w_0_0# gnd 0.10fF
C423 ffi_0/nand_6/a ffi_0/inv_1/op 0.13fF
C424 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C425 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C426 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_1/b 0.31fF
C427 sumffo_1/ffo_0/d ffi_0/q 0.27fF
C428 gnd ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C429 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C430 cla_0/g0 ffi_0/q 0.08fF
C431 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/inv_1/w_0_6# 0.04fF
C432 gnd z2o 0.80fF
C433 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C434 ffipg_2/ffi_0/nand_2/w_0_0# ffipg_2/ffi_0/nand_3/a 0.04fF
C435 ffipg_1/ffi_0/nand_2/w_0_0# gnd 0.10fF
C436 sumffo_3/ffo_0/inv_0/w_0_6# gnd 0.07fF
C437 sumffo_1/ffo_0/nand_2/w_0_0# gnd 0.10fF
C438 clk sumffo_1/ffo_0/nand_3/b 0.33fF
C439 gnd nand_2/b 1.90fF
C440 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# 0.04fF
C441 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C442 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q 0.32fF
C443 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b 0.13fF
C444 sumffo_0/ffo_0/inv_1/w_0_6# gnd 0.06fF
C445 ffipg_3/ffi_0/nand_1/a clk 0.13fF
C446 gnd ffipg_0/ffi_0/nand_3/w_0_0# 0.11fF
C447 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C448 ffo_0/nand_3/a gnd 0.49fF
C449 inv_5/in gnd 0.49fF
C450 ffo_0/inv_0/op gnd 0.37fF
C451 inv_5/w_0_6# cla_0/n 0.06fF
C452 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C453 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a 0.31fF
C454 clk ffipg_0/ffi_1/nand_3/a 0.13fF
C455 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C456 clk sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C457 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C458 ffi_0/nand_2/w_0_0# ffi_0/nand_3/a 0.04fF
C459 gnd ffipg_3/ffi_1/nand_7/w_0_0# 0.10fF
C460 sumffo_2/xor_0/a_10_10# gnd 0.93fF
C461 clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C462 cla_0/l cla_2/p1 0.30fF
C463 cla_2/p1 cla_2/nor_0/w_0_0# 0.06fF
C464 ffipg_3/pggen_0/xor_0/a_10_10# gnd 0.93fF
C465 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k 0.52fF
C466 ffipg_2/ffi_0/nand_3/b gnd 0.74fF
C467 gnd ffipg_1/ffi_0/nand_6/a 0.37fF
C468 ffipg_0/ffi_0/q ffipg_0/k 0.07fF
C469 ffi_0/nand_6/a ffi_0/q 0.31fF
C470 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/inv_1/op 0.33fF
C471 sumffo_1/xor_0/inv_1/op nand_2/b 0.22fF
C472 ffi_0/nand_3/b ffi_0/nand_3/a 0.31fF
C473 gnd ffipg_0/ffi_1/nand_3/b 0.74fF
C474 cla_1/l nand_2/b 0.31fF
C475 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C476 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C477 ffipg_1/ffi_0/nand_1/a gnd 0.44fF
C478 nor_1/b inv_1/in 0.16fF
C479 inv_1/op sumffo_2/xor_0/inv_0/op 0.27fF
C480 sumffo_2/ffo_0/nand_0/b gnd 0.63fF
C481 cla_0/l cla_2/inv_0/in 0.16fF
C482 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/w_0_0# 0.04fF
C483 nor_0/w_0_0# nor_0/b 0.06fF
C484 sumffo_1/ffo_0/nand_4/w_0_0# gnd 0.10fF
C485 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# 0.04fF
C486 gnd ffipg_1/ffi_0/nand_0/a_13_n26# 0.01fF
C487 gnd ffi_0/nand_1/a 0.44fF
C488 nor_1/w_0_0# cla_0/n 0.06fF
C489 inv_1/in gnd 0.33fF
C490 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C491 ffipg_0/k ffi_0/q 0.19fF
C492 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a 0.00fF
C493 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/qbar 0.06fF
C494 cla_1/p0 cla_0/g0 0.38fF
C495 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_6/a 0.04fF
C496 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b 0.32fF
C497 x4in ffipg_3/ffi_1/inv_1/op 0.01fF
C498 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C499 clk sumffo_0/ffo_0/nand_0/b 0.04fF
C500 ffipg_2/ffi_0/q ffipg_2/ffi_1/q 0.73fF
C501 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C502 ffipg_3/k ffipg_3/ffi_0/q 0.07fF
C503 ffipg_2/ffi_0/nand_4/w_0_0# gnd 0.10fF
C504 ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C505 gnd ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C506 clk ffipg_3/ffi_1/inv_1/op 0.07fF
C507 ffipg_2/ffi_1/nand_1/b gnd 0.57fF
C508 ffipg_0/pggen_0/nor_0/w_0_0# gnd 0.11fF
C509 sumffo_0/ffo_0/nand_6/w_0_0# gnd 0.10fF
C510 clk y3in 0.68fF
C511 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C512 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# 0.04fF
C513 ffo_0/nand_6/a clk 0.13fF
C514 sumffo_3/ffo_0/nand_0/w_0_0# gnd 0.10fF
C515 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C516 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# 0.04fF
C517 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C518 sumffo_1/ffo_0/inv_1/w_0_6# gnd 0.06fF
C519 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_1/b 0.04fF
C520 ffipg_0/ffi_1/nand_7/w_0_0# gnd 0.10fF
C521 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_3/b 0.04fF
C522 gnd ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C523 gnd ffipg_3/ffi_1/q 2.24fF
C524 nor_0/w_0_0# inv_0/in 0.11fF
C525 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C526 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar 0.32fF
C527 ffipg_1/ffi_1/inv_0/op x2in 0.04fF
C528 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C529 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/q 0.00fF
C530 sumffo_1/xor_0/inv_0/w_0_6# gnd 0.09fF
C531 sumffo_3/ffo_0/nand_3/w_0_0# gnd 0.11fF
C532 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C533 nor_0/w_0_0# gnd 0.46fF
C534 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C535 clk ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C536 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C537 ffipg_2/ffi_1/nand_6/w_0_0# gnd 0.10fF
C538 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b 0.13fF
C539 gnd ffipg_2/ffi_1/nand_0/a_13_n26# 0.01fF
C540 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_0/op 0.32fF
C541 ffipg_1/ffi_0/q ffipg_1/ffi_1/q 0.73fF
C542 cla_2/p1 gnd 1.00fF
C543 ffipg_2/ffi_0/nand_1/a gnd 0.44fF
C544 gnd ffipg_1/ffi_0/inv_1/op 1.85fF
C545 ffipg_0/ffi_1/inv_0/op ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C546 clk ffo_0/nand_0/b 0.04fF
C547 sumffo_3/xor_0/a_10_10# ffi_0/q 0.04fF
C548 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_3/b 0.00fF
C549 ffipg_1/ffi_1/nand_7/w_0_0# gnd 0.10fF
C550 sumffo_2/ffo_0/inv_0/op gnd 0.51fF
C551 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C552 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_3/b 0.04fF
C553 cla_2/inv_0/in gnd 0.34fF
C554 clk sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C555 nor_0/w_0_0# inv_0/op 0.10fF
C556 gnd ffipg_3/ffi_1/inv_0/op 0.27fF
C557 ffipg_2/ffi_0/nand_3/a gnd 0.33fF
C558 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/inv_1/op 0.33fF
C559 sumffo_1/ffo_0/nand_3/w_0_0# gnd 0.11fF
C560 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_3/b 0.00fF
C561 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C562 sumffo_3/xor_0/inv_1/op ffipg_3/k 0.22fF
C563 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C564 clk ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C565 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/b 0.31fF
C566 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q 0.27fF
C567 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C568 inv_1/in inv_1/op 0.04fF
C569 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C570 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C571 ffipg_1/ffi_1/nand_1/a gnd 0.44fF
C572 nor_2/w_0_0# gnd 0.15fF
C573 sumffo_0/ffo_0/nand_7/a gnd 0.33fF
C574 inv_5/w_0_6# cla_2/l 0.08fF
C575 gnd couto 0.80fF
C576 sumffo_3/ffo_0/nand_1/b gnd 0.57fF
C577 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/q 0.00fF
C578 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C579 ffipg_0/ffi_0/nand_0/w_0_0# gnd 0.10fF
C580 nor_3/w_0_0# cla_2/n 0.06fF
C581 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C582 gnd ffi_0/inv_0/op 0.27fF
C583 ffipg_1/ffi_0/inv_0/op ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C584 sumffo_1/xor_0/w_n3_4# sumffo_1/ffo_0/d 0.02fF
C585 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/d 0.40fF
C586 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# 0.04fF
C587 cla_1/n inv_4/in 0.02fF
C588 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C589 gnd sumffo_3/ffo_0/nand_7/a 0.33fF
C590 ffi_0/nand_7/a ffi_0/q 0.00fF
C591 ffipg_2/ffi_1/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C592 ffipg_1/ffi_1/nand_5/w_0_0# gnd 0.10fF
C593 gnd y1in 0.22fF
C594 nor_4/b nor_3/w_0_0# 0.03fF
C595 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C596 y3in ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C597 gnd ffo_0/nand_6/w_0_0# 0.10fF
C598 clk ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C599 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/nand_1/a 0.04fF
C600 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C601 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.35fF
C602 gnd ffipg_1/ffi_1/nand_2/w_0_0# 0.10fF
C603 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# 0.04fF
C604 clk ffipg_0/ffi_0/inv_1/op 0.07fF
C605 gnd ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C606 ffipg_2/ffi_1/nand_0/w_0_0# ffipg_2/ffi_1/nand_1/a 0.04fF
C607 cla_0/l ffipg_2/ffi_0/q 0.13fF
C608 clk x2in 0.68fF
C609 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C610 clk ffo_0/nand_3/b 0.33fF
C611 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/d 0.06fF
C612 ffipg_3/ffi_1/nand_6/a gnd 0.37fF
C613 ffipg_3/ffi_1/inv_0/w_0_6# gnd 0.06fF
C614 ffipg_1/ffi_1/inv_1/w_0_6# gnd 0.06fF
C615 ffipg_0/ffi_1/nand_2/w_0_0# gnd 0.10fF
C616 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_1/w_0_6# 0.03fF
C617 gnd sumffo_1/ffo_0/nand_5/w_0_0# 0.10fF
C618 cla_0/l inv_2/w_0_6# 0.06fF
C619 ffipg_1/ffi_1/inv_0/w_0_6# gnd 0.06fF
C620 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C621 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_7/a 0.04fF
C622 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/b 0.31fF
C623 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C624 cla_0/l ffi_0/q 0.33fF
C625 ffo_0/nand_7/a couto 0.00fF
C626 cla_0/l cla_2/g1 0.26fF
C627 nor_2/b inv_3/w_0_6# 0.03fF
C628 ffipg_2/ffi_1/nand_3/b gnd 0.74fF
C629 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C630 ffipg_3/ffi_0/qbar gnd 0.67fF
C631 clk ffipg_0/ffi_0/nand_2/w_0_0# 0.06fF
C632 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C633 sumffo_0/ffo_0/nand_0/a_13_n26# gnd 0.01fF
C634 gnd ffipg_3/ffi_0/nand_1/w_0_0# 0.10fF
C635 ffo_0/nand_3/w_0_0# ffo_0/nand_3/b 0.06fF
C636 ffipg_2/ffi_1/qbar gnd 0.67fF
C637 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/qbar 0.00fF
C638 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/d 0.06fF
C639 ffipg_0/ffi_0/inv_0/op clk 0.32fF
C640 cla_0/inv_0/in cla_0/inv_0/op 0.04fF
C641 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b 0.13fF
C642 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a 0.31fF
C643 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/inv_1/op 0.13fF
C644 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C645 nor_0/w_0_0# nand_2/b 0.04fF
C646 sumffo_2/ffo_0/nand_4/w_0_0# clk 0.06fF
C647 sumffo_3/ffo_0/d ffi_0/q 0.16fF
C648 nor_0/b ffi_0/q 0.32fF
C649 nor_3/b nor_3/w_0_0# 0.06fF
C650 ffo_0/qbar gnd 0.62fF
C651 sumffo_2/ffo_0/nand_1/b gnd 0.57fF
C652 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/w_0_0# 0.06fF
C653 clk cinin 0.68fF
C654 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C655 ffipg_2/ffi_0/nand_3/w_0_0# gnd 0.11fF
C656 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q 0.27fF
C657 clk ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C658 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_4/w_0_0# 0.04fF
C659 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C660 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C661 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C662 inv_2/in inv_2/w_0_6# 0.10fF
C663 ffi_0/inv_1/op gnd 1.89fF
C664 clk sumffo_0/ffo_0/nand_1/b 0.45fF
C665 sumffo_2/ffo_0/nand_6/w_0_0# gnd 0.10fF
C666 ffipg_3/ffi_0/nand_0/w_0_0# gnd 0.10fF
C667 ffipg_2/ffi_0/inv_0/op gnd 0.27fF
C668 gnd sumffo_1/ffo_0/nand_1/a 0.44fF
C669 inv_2/in ffi_0/q 0.13fF
C670 cla_0/inv_0/in cla_0/g0 0.16fF
C671 ffipg_3/ffi_0/nand_2/w_0_0# y4in 0.06fF
C672 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C673 sumffo_3/ffo_0/nand_2/w_0_0# gnd 0.10fF
C674 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/sbar 0.06fF
C675 clk ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C676 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_1/b 0.45fF
C677 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/ffo_0/nand_7/a 0.06fF
C678 z3o sumffo_2/ffo_0/nand_7/a 0.00fF
C679 clk ffipg_0/ffi_0/nand_1/a 0.13fF
C680 ffipg_0/ffi_1/q ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C681 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b 0.13fF
C682 ffo_0/nand_5/w_0_0# gnd 0.10fF
C683 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C684 clk ffi_0/nand_2/w_0_0# 0.06fF
C685 sumffo_0/ffo_0/nand_3/b gnd 0.74fF
C686 ffipg_0/ffi_0/nand_7/a gnd 0.37fF
C687 ffipg_0/pggen_0/xor_0/inv_1/op gnd 0.35fF
C688 inv_6/in gnd 0.33fF
C689 sumffo_1/sbar sumffo_1/ffo_0/nand_7/a 0.31fF
C690 ffipg_0/ffi_0/q gnd 3.00fF
C691 y2in ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C692 ffipg_0/ffi_1/q ffipg_0/k 0.46fF
C693 clk sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C694 sumffo_0/ffo_0/nand_2/w_0_0# gnd 0.10fF
C695 ffipg_1/k ffi_0/q 0.06fF
C696 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C697 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a 0.13fF
C698 sumffo_0/xor_0/inv_1/op ffi_0/q 0.22fF
C699 cla_0/l cla_1/p0 0.09fF
C700 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a 0.00fF
C701 nor_1/b inv_2/w_0_6# 0.03fF
C702 inv_0/in ffi_0/q 0.07fF
C703 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_3/b 0.00fF
C704 ffipg_2/ffi_0/q gnd 3.00fF
C705 gnd ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C706 ffipg_0/ffi_0/inv_0/w_0_6# gnd 0.06fF
C707 ffo_0/nand_7/a ffo_0/qbar 0.31fF
C708 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/nand_3/a 0.04fF
C709 cla_0/n ffipg_3/k 0.06fF
C710 ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_3/b 0.31fF
C711 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C712 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a 0.13fF
C713 gnd inv_2/w_0_6# 0.17fF
C714 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C715 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a 0.31fF
C716 nor_3/b cla_2/n 0.41fF
C717 gnd ffo_0/nand_1/b 0.57fF
C718 cla_2/p0 ffipg_3/k 0.06fF
C719 nor_2/b gnd 0.32fF
C720 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_0/op 0.32fF
C721 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C722 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# 0.04fF
C723 sumffo_0/xor_0/inv_1/w_0_6# ffi_0/q 0.23fF
C724 gnd ffi_0/q 2.14fF
C725 clk ffipg_1/ffi_1/inv_1/op 0.07fF
C726 cla_2/g1 gnd 0.65fF
C727 inv_8/w_0_6# ffi_0/q 0.06fF
C728 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/k 0.01fF
C729 inv_4/op gnd 0.58fF
C730 ffo_0/nand_0/w_0_0# ffo_0/nand_0/b 0.06fF
C731 cla_0/g0 nor_0/a 0.68fF
C732 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_3/b 0.31fF
C733 inv_7/op inv_7/w_0_6# 0.03fF
C734 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C735 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_3/b 0.33fF
C736 ffi_0/nand_3/b ffi_0/nand_4/w_0_0# 0.06fF
C737 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k 0.06fF
C738 ffo_0/nand_7/a ffo_0/nand_5/w_0_0# 0.04fF
C739 sumffo_2/ffo_0/d gnd 0.41fF
C740 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/nand_7/a 0.06fF
C741 ffipg_1/ffi_1/nand_3/a gnd 0.33fF
C742 ffo_0/nand_7/w_0_0# gnd 0.10fF
C743 ffipg_1/ffi_0/inv_0/op gnd 0.27fF
C744 gnd ffipg_1/ffi_0/nand_1/b 0.57fF
C745 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q 0.22fF
C746 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C747 ffo_0/nand_0/b ffo_0/d 0.40fF
C748 cla_0/nor_0/w_0_0# gnd 0.31fF
C749 clk ffi_0/nand_0/w_0_0# 0.06fF
C750 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/nand_6/a 0.06fF
C751 ffipg_0/ffi_1/nand_0/w_0_0# ffipg_0/ffi_1/inv_0/op 0.06fF
C752 ffipg_3/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C753 ffipg_3/ffi_0/nand_6/a gnd 0.37fF
C754 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C755 clk sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C756 sumffo_1/xor_0/inv_1/op ffi_0/q 0.04fF
C757 cla_2/p1 ffipg_3/ffi_1/q 0.22fF
C758 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b 0.32fF
C759 cla_0/nor_1/w_0_0# cla_0/g0 0.06fF
C760 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C761 gnd ffipg_3/ffi_1/qbar 0.67fF
C762 ffo_0/nand_7/a ffo_0/nand_1/b 0.13fF
C763 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/b 0.31fF
C764 gnd ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C765 cla_1/p0 ffipg_1/k 0.05fF
C766 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_3/a 0.04fF
C767 sumffo_3/xor_0/w_n3_4# ffi_0/q 0.01fF
C768 ffipg_3/ffi_1/nand_2/w_0_0# ffipg_3/ffi_1/nand_3/a 0.04fF
C769 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C770 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar 0.32fF
C771 clk ffipg_0/ffi_0/nand_3/a 0.13fF
C772 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C773 ffo_0/nand_0/b ffo_0/nand_2/w_0_0# 0.06fF
C774 gnd sumffo_1/ffo_0/nand_1/w_0_0# 0.10fF
C775 sumffo_0/ffo_0/inv_0/w_0_6# sumffo_0/ffo_0/d 0.06fF
C776 gnd z1o 0.80fF
C777 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/qbar 0.31fF
C778 sumffo_3/xor_0/w_n3_4# inv_4/op 0.06fF
C779 sumffo_0/ffo_0/nand_6/a z1o 0.31fF
C780 sumffo_2/xor_0/inv_0/op ffi_0/q 0.06fF
C781 gnd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C782 gnd ffipg_0/ffi_1/nand_1/b 0.57fF
C783 ffo_0/nand_7/a ffo_0/nand_7/w_0_0# 0.06fF
C784 cla_1/p0 gnd 1.06fF
C785 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/inv_1/op 0.45fF
C786 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a 0.00fF
C787 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C788 sumffo_3/ffo_0/nand_6/a clk 0.13fF
C789 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_7/a 0.04fF
C790 ffipg_1/ffi_0/nand_3/a gnd 0.33fF
C791 cla_2/p1 cla_2/inv_0/in 0.02fF
C792 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b 0.32fF
C793 sumffo_2/ffo_0/nand_3/a gnd 0.33fF
C794 gnd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C795 ffo_0/d ffo_0/nand_2/w_0_0# 0.06fF
C796 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op 0.06fF
C797 ffipg_2/ffi_1/nand_7/a gnd 0.37fF
C798 nor_0/a ffipg_0/k 0.05fF
C799 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C800 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C801 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C802 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C803 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C804 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_3/b 0.00fF
C805 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/b 0.31fF
C806 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# 0.04fF
C807 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/qbar 0.06fF
C808 gnd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C809 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C810 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C811 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_3/b 0.06fF
C812 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C813 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/a 0.06fF
C814 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_1/w_0_6# 0.03fF
C815 clk sumffo_1/ffo_0/d 0.04fF
C816 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_1/q 0.06fF
C817 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C818 ffipg_3/ffi_0/inv_1/op gnd 1.85fF
C819 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C820 nand_2/b inv_2/w_0_6# 0.03fF
C821 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C822 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b 0.32fF
C823 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C824 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C825 cla_1/l cla_1/p0 0.16fF
C826 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/q 0.31fF
C827 gnd ffipg_2/ffi_0/nand_7/a 0.37fF
C828 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C829 nand_2/b ffi_0/q 0.04fF
C830 ffi_0/nand_7/w_0_0# ffi_0/nand_7/a 0.06fF
C831 ffipg_0/ffi_1/nand_3/w_0_0# gnd 0.11fF
C832 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/inv_1/op 0.45fF
C833 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C834 inv_9/in nor_4/a 0.02fF
C835 sumffo_1/ffo_0/nand_2/a_13_n26# gnd 0.01fF
C836 sumffo_3/sbar z4o 0.32fF
C837 ffipg_2/ffi_1/nand_7/w_0_0# ffipg_2/ffi_1/q 0.04fF
C838 sumffo_0/xor_0/w_n3_4# gnd 0.12fF
C839 y2in gnd 0.22fF
C840 gnd y4in 0.22fF
C841 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C842 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C843 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C844 sumffo_3/ffo_0/nand_4/w_0_0# gnd 0.10fF
C845 ffipg_3/ffi_1/inv_1/w_0_6# clk 0.06fF
C846 clk ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C847 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op 0.06fF
C848 gnd sumffo_2/xor_0/inv_1/op 0.35fF
C849 sumffo_0/ffo_0/inv_0/w_0_6# sumffo_0/ffo_0/inv_0/op 0.03fF
C850 sumffo_2/xor_0/a_10_10# ffi_0/q 0.04fF
C851 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C852 ffipg_0/ffi_1/inv_0/op x1in 0.04fF
C853 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_1/b 0.04fF
C854 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C855 ffipg_3/ffi_0/inv_0/op gnd 0.27fF
C856 ffipg_3/ffi_1/inv_0/w_0_6# ffipg_3/ffi_1/inv_0/op 0.03fF
C857 gnd ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C858 ffi_0/inv_0/w_0_6# gnd 0.06fF
C859 ffipg_2/pggen_0/xor_0/inv_0/op gnd 0.32fF
C860 gnd ffo_0/inv_0/w_0_6# 0.07fF
C861 sumffo_1/xor_0/w_n3_4# ffipg_1/k 0.06fF
C862 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/qbar 0.04fF
C863 ffo_0/nand_6/w_0_0# couto 0.06fF
C864 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a 0.13fF
C865 sumffo_2/xor_0/a_10_10# sumffo_2/ffo_0/d 0.45fF
C866 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C867 gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C868 nor_4/a nor_4/w_0_0# 0.07fF
C869 clk ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C870 ffipg_2/pggen_0/nor_0/w_0_0# cla_2/p0 0.05fF
C871 ffipg_0/ffi_0/q ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C872 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C873 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# 0.04fF
C874 gnd ffi_0/nand_3/a 0.33fF
C875 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C876 ffipg_0/ffi_0/inv_1/w_0_6# ffipg_0/ffi_0/inv_1/op 0.04fF
C877 ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_3/b 0.31fF
C878 cla_2/l inv_7/w_0_6# 0.06fF
C879 cla_0/l cla_0/inv_0/in 0.07fF
C880 ffipg_1/ffi_1/q ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C881 sumffo_0/ffo_0/d gnd 0.41fF
C882 ffi_0/nand_1/b ffi_0/nand_1/w_0_0# 0.06fF
C883 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C884 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/d 0.40fF
C885 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C886 ffipg_0/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C887 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/inv_1/op 0.33fF
C888 ffi_0/nand_7/w_0_0# nor_0/b 0.06fF
C889 ffi_0/nand_4/w_0_0# ffi_0/nand_6/a 0.04fF
C890 inv_9/in gnd 0.33fF
C891 sumffo_1/xor_0/w_n3_4# gnd 0.12fF
C892 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C893 sumffo_1/ffo_0/nand_0/b gnd 0.62fF
C894 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar 0.32fF
C895 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/q 0.31fF
C896 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# 0.04fF
C897 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_1/b 0.31fF
C898 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C899 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C900 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C901 ffipg_1/ffi_0/nand_2/w_0_0# ffipg_1/ffi_0/nand_3/a 0.04fF
C902 ffipg_0/ffi_1/nand_0/w_0_0# gnd 0.10fF
C903 ffipg_3/ffi_1/nand_7/w_0_0# ffipg_3/ffi_1/qbar 0.06fF
C904 gnd ffipg_2/ffi_0/qbar 0.67fF
C905 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C906 ffi_0/nand_1/b ffi_0/nand_3/w_0_0# 0.04fF
C907 clk ffipg_3/ffi_1/nand_3/a 0.13fF
C908 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/ffi_1/q 0.06fF
C909 clk ffipg_2/ffi_1/inv_0/op 0.32fF
C910 ffipg_0/ffi_1/inv_1/op x1in 0.01fF
C911 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C912 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_3/a 0.06fF
C913 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C914 cla_2/nor_1/w_0_0# gnd 0.31fF
C915 gnd ffipg_1/ffi_1/nand_6/w_0_0# 0.10fF
C916 gnd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C917 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_3/b 0.06fF
C918 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a 0.31fF
C919 gnd ffo_0/nand_4/w_0_0# 0.10fF
C920 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_0/op 0.08fF
C921 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_1/q 0.06fF
C922 gnd ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C923 ffo_0/qbar couto 0.32fF
C924 sumffo_3/xor_0/inv_0/w_0_6# gnd 0.09fF
C925 ffipg_2/k cla_0/n 0.06fF
C926 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/qbar 0.04fF
C927 ffipg_1/ffi_0/nand_4/w_0_0# gnd 0.10fF
C928 ffipg_0/ffi_1/q gnd 2.24fF
C929 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/k 0.21fF
C930 gnd sumffo_0/sbar 0.62fF
C931 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C932 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_1/a 0.04fF
C933 ffipg_2/k cla_2/p0 0.05fF
C934 gnd nor_4/w_0_0# 0.15fF
C935 sumffo_0/ffo_0/nand_6/a sumffo_0/sbar 0.00fF
C936 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/w_0_0# 0.04fF
C937 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/w_0_0# 0.04fF
C938 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C939 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C940 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b 0.32fF
C941 inv_5/w_0_6# gnd 0.41fF
C942 nor_0/w_0_0# ffi_0/q 0.16fF
C943 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C944 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C945 ffipg_1/ffi_1/q ffipg_1/k 0.46fF
C946 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C947 cla_0/l nor_0/a 0.16fF
C948 ffipg_1/ffi_1/inv_1/op x2in 0.01fF
C949 sumffo_0/ffo_0/nand_3/w_0_0# gnd 0.11fF
C950 ffo_0/qbar ffo_0/nand_6/w_0_0# 0.04fF
C951 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_3/b 0.04fF
C952 clk ffo_0/inv_1/w_0_6# 0.06fF
C953 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C954 ffipg_1/ffi_0/qbar gnd 0.67fF
C955 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C956 ffipg_3/ffi_0/nand_2/w_0_0# clk 0.06fF
C957 ffi_0/nand_3/b ffi_0/nand_1/w_0_0# 0.04fF
C958 clk ffipg_2/ffi_1/inv_1/op 0.07fF
C959 ffipg_1/ffi_0/nand_2/w_0_0# y2in 0.06fF
C960 cla_2/g1 cla_2/p1 0.00fF
C961 ffi_0/nand_7/w_0_0# gnd 0.10fF
C962 clk sumffo_2/ffo_0/nand_3/b 0.33fF
C963 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/ffi_1/q 0.06fF
C964 sumffo_2/ffo_0/nand_6/a gnd 0.33fF
C965 ffipg_0/ffi_0/nand_7/w_0_0# ffipg_0/ffi_0/qbar 0.06fF
C966 ffipg_3/pggen_0/nor_0/w_0_0# gnd 0.11fF
C967 ffi_0/nand_2/w_0_0# cinin 0.06fF
C968 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.32fF
C969 sumffo_0/ffo_0/nand_6/w_0_0# z1o 0.06fF
C970 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C971 nor_3/b cla_2/l 0.10fF
C972 ffi_0/nand_3/b ffi_0/nand_3/w_0_0# 0.06fF
C973 ffi_0/nand_3/b ffi_0/nand_1/b 0.32fF
C974 ffipg_1/ffi_1/q gnd 2.24fF
C975 nor_1/w_0_0# nor_1/b 0.06fF
C976 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/ffo_0/nand_6/a 0.06fF
C977 cla_2/g1 cla_2/inv_0/in 0.04fF
C978 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C979 ffipg_3/ffi_1/inv_1/w_0_6# ffipg_3/ffi_1/inv_1/op 0.04fF
C980 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar 0.32fF
C981 ffipg_0/pggen_0/xor_0/inv_0/op gnd 0.32fF
C982 nor_0/b nor_0/a 0.32fF
C983 clk ffipg_0/ffi_1/inv_0/op 0.32fF
C984 sumffo_0/ffo_0/inv_0/op gnd 0.27fF
C985 ffipg_2/ffi_0/nand_2/w_0_0# clk 0.06fF
C986 nor_1/w_0_0# gnd 0.15fF
C987 cla_0/inv_0/in gnd 0.34fF
C988 nor_2/w_0_0# nor_2/b 0.06fF
C989 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_1/b 0.45fF
C990 sumffo_3/ffo_0/nand_6/a sumffo_3/sbar 0.00fF
C991 gnd ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C992 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d 0.04fF
C993 sumffo_1/ffo_0/nand_6/a gnd 0.33fF
C994 sumffo_2/ffo_0/nand_7/a sumffo_2/sbar 0.31fF
C995 ffipg_3/ffi_1/nand_2/w_0_0# gnd 0.10fF
C996 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_1/b 0.13fF
C997 clk x3in 0.68fF
C998 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_3/b 0.06fF
C999 ffipg_0/ffi_0/inv_0/w_0_6# y1in 0.06fF
C1000 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b 0.32fF
C1001 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C1002 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a 0.00fF
C1003 nor_2/w_0_0# inv_4/op 0.03fF
C1004 ffipg_0/ffi_0/nand_1/w_0_0# ffipg_0/ffi_0/nand_3/b 0.04fF
C1005 gnd sumffo_1/xor_0/a_10_10# 0.93fF
C1006 sumffo_1/ffo_0/nand_1/b gnd 0.57fF
C1007 ffi_0/nand_1/b ffi_0/nand_5/w_0_0# 0.06fF
C1008 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C1009 ffipg_2/ffi_0/inv_1/w_0_6# ffipg_2/ffi_0/inv_1/op 0.04fF
C1010 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# 0.04fF
C1011 ffo_0/inv_0/op ffo_0/inv_0/w_0_6# 0.03fF
C1012 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_0/b 0.06fF
C1013 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C1014 ffo_0/nand_7/w_0_0# couto 0.04fF
C1015 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C1016 inv_3/in inv_3/w_0_6# 0.10fF
C1017 nor_0/a ffipg_1/k 0.06fF
C1018 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/xor_0/inv_0/op 0.03fF
C1019 cla_2/l cla_0/n 0.32fF
C1020 ffipg_2/k sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C1021 ffipg_1/ffi_1/nand_3/w_0_0# ffipg_1/ffi_1/nand_3/b 0.06fF
C1022 gnd x1in 0.22fF
C1023 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/d 0.40fF
C1024 ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_2/w_0_0# 0.04fF
C1025 cla_2/p0 cla_2/l 0.16fF
C1026 cla_2/nand_0/a_13_n26# gnd 0.01fF
C1027 nor_0/a inv_0/in 0.02fF
C1028 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/w_0_0# 0.06fF
C1029 clk ffipg_2/ffi_0/inv_1/op 0.07fF
C1030 clk ffipg_0/ffi_1/inv_1/op 0.07fF
C1031 gnd ffipg_1/ffi_1/nand_3/w_0_0# 0.11fF
C1032 gnd ffipg_3/ffi_1/nand_6/w_0_0# 0.10fF
C1033 clk ffipg_3/ffi_0/nand_3/a 0.13fF
C1034 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op 0.13fF
C1035 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1036 nor_0/a gnd 0.54fF
C1037 sumffo_0/ffo_0/nand_7/a z1o 0.00fF
C1038 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# 0.04fF
C1039 cla_0/l cla_0/nand_0/w_0_0# 0.06fF
C1040 sumffo_3/xor_0/a_10_10# ffipg_3/k 0.12fF
C1041 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C1042 ffipg_1/ffi_1/inv_0/op gnd 0.27fF
C1043 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_3/a 0.06fF
C1044 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C1045 gnd ffi_0/inv_1/w_0_6# 0.06fF
C1046 sumffo_0/ffo_0/nand_0/w_0_0# gnd 0.10fF
C1047 gnd ffipg_3/ffi_1/nand_0/w_0_0# 0.10fF
C1048 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C1049 gnd sumffo_2/ffo_0/nand_7/a 0.33fF
C1050 ffipg_2/ffi_1/nand_7/w_0_0# gnd 0.10fF
C1051 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C1052 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C1053 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C1054 cla_0/nor_1/w_0_0# gnd 0.31fF
C1055 sumffo_2/xor_0/a_38_n43# ffi_0/q 0.01fF
C1056 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# 0.16fF
C1057 inv_5/in inv_5/w_0_6# 0.10fF
C1058 clk sumffo_3/ffo_0/d 0.04fF
C1059 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1060 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/qbar 0.00fF
C1061 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C1062 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a 0.00fF
C1063 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C1064 nor_1/w_0_0# inv_1/op 0.03fF
C1065 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C1066 clk nor_4/a 0.03fF
C1067 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/nand_6/a 0.04fF
C1068 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/qbar 0.00fF
C1069 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/inv_0/op 0.06fF
C1070 sumffo_3/ffo_0/nand_0/b gnd 0.53fF
C1071 gnd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C1072 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C1073 ffipg_3/ffi_1/nand_0/w_0_0# ffipg_3/ffi_1/nand_1/a 0.04fF
C1074 y2in ffipg_1/ffi_0/inv_1/op 0.01fF
C1075 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1076 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C1077 sumffo_1/ffo_0/nand_6/a z2o 0.31fF
C1078 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C1079 inv_3/in gnd 0.47fF
C1080 ffipg_3/ffi_0/nand_7/w_0_0# gnd 0.10fF
C1081 gnd inv_4/in 0.33fF
C1082 ffipg_2/ffi_0/nand_2/w_0_0# y3in 0.06fF
C1083 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a 0.00fF
C1084 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/inv_1/op 0.45fF
C1085 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C1086 cla_0/inv_0/w_0_6# cla_0/inv_0/op 0.03fF
C1087 gnd sumffo_1/ffo_0/nand_3/a 0.48fF
C1088 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/nand_7/a 0.06fF
C1089 ffipg_2/ffi_0/inv_1/w_0_6# gnd 0.06fF
C1090 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/b 0.31fF
C1091 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C1092 ffipg_2/ffi_1/inv_1/w_0_6# ffipg_2/ffi_1/inv_1/op 0.04fF
C1093 cla_0/l ffipg_3/k 0.10fF
C1094 gnd x4in 0.22fF
C1095 inv_2/w_0_6# ffi_0/q 0.06fF
C1096 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b 0.32fF
C1097 gnd ffipg_0/ffi_1/nand_1/a 0.45fF
C1098 ffo_0/nand_0/b ffo_0/inv_1/w_0_6# 0.03fF
C1099 sumffo_3/ffo_0/nand_1/a gnd 0.33fF
C1100 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1101 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/ffi_1/q 0.06fF
C1102 sumffo_2/ffo_0/nand_1/w_0_0# gnd 0.10fF
C1103 ffipg_2/ffi_0/inv_0/op ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C1104 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/sbar 0.04fF
C1105 clk gnd 24.51fF
C1106 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C1107 clk sumffo_0/ffo_0/nand_6/a 0.13fF
C1108 cla_0/nand_0/w_0_0# gnd 0.10fF
C1109 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/qbar 0.31fF
C1110 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C1111 gnd ffipg_2/ffi_1/nand_1/a 0.44fF
C1112 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/q 0.04fF
C1113 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C1114 ffipg_2/ffi_1/nand_4/w_0_0# ffipg_2/ffi_1/inv_1/op 0.06fF
C1115 ffipg_2/ffi_0/nand_6/a gnd 0.37fF
C1116 ffipg_2/pggen_0/xor_0/inv_1/op gnd 0.35fF
C1117 sumffo_2/ffo_0/d ffi_0/q 0.27fF
C1118 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/nand_7/a 0.04fF
C1119 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C1120 y3in ffipg_2/ffi_0/inv_1/op 0.01fF
C1121 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k 0.52fF
C1122 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C1123 nor_1/w_0_0# inv_1/in 0.11fF
C1124 ffi_0/inv_0/w_0_6# ffi_0/inv_0/op 0.03fF
C1125 sumffo_1/sbar gnd 0.62fF
C1126 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C1127 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_6/a 0.04fF
C1128 cla_1/nor_1/w_0_0# gnd 0.31fF
C1129 ffi_0/nand_4/w_0_0# gnd 0.10fF
C1130 ffo_0/nand_3/w_0_0# gnd 0.11fF
C1131 ffo_0/nand_1/a ffo_0/nand_0/b 0.13fF
C1132 cla_0/l inv_7/w_0_6# 0.06fF
C1133 ffipg_1/ffi_1/nand_0/w_0_0# clk 0.06fF
C1134 gnd ffipg_3/ffi_0/q 3.00fF
C1135 clk ffipg_3/ffi_1/nand_1/a 0.13fF
C1136 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/ffi_1/q 0.06fF
C1137 ffipg_3/ffi_1/nand_4/w_0_0# gnd 0.10fF
C1138 ffipg_1/pggen_0/xor_0/inv_1/op gnd 0.35fF
C1139 gnd sumffo_1/xor_0/inv_0/op 0.32fF
C1140 gnd sumffo_1/ffo_0/nand_3/b 0.74fF
C1141 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C1142 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/q 0.31fF
C1143 cla_2/p0 ffipg_2/ffi_1/q 0.22fF
C1144 ffipg_0/ffi_0/nand_6/a gnd 0.37fF
C1145 ffo_0/nand_1/a ffo_0/nand_0/w_0_0# 0.04fF
C1146 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C1147 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/b 0.31fF
C1148 sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d 0.52fF
C1149 sumffo_2/ffo_0/nand_3/w_0_0# gnd 0.11fF
C1150 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/q 0.00fF
C1151 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_1/q 0.06fF
C1152 ffipg_1/ffi_0/nand_5/w_0_0# gnd 0.10fF
C1153 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1154 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/ffi_1/q 0.06fF
C1155 ffipg_3/ffi_0/nand_1/a gnd 0.44fF
C1156 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C1157 sumffo_1/ffo_0/nand_6/w_0_0# z2o 0.06fF
C1158 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C1159 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b 0.32fF
C1160 ffipg_0/ffi_1/nand_3/a gnd 0.33fF
C1161 sumffo_2/ffo_0/inv_1/w_0_6# gnd 0.07fF
C1162 cla_1/inv_0/op cla_0/n 0.02fF
C1163 ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C1164 ffipg_1/ffi_1/nand_1/b gnd 0.57fF
C1165 sumffo_0/ffo_0/nand_7/a sumffo_0/sbar 0.31fF
C1166 sumffo_0/ffo_0/nand_4/w_0_0# gnd 0.10fF
C1167 nor_3/w_0_0# gnd 0.15fF
C1168 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# 0.04fF
C1169 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C1170 ffipg_2/ffi_1/nand_3/a clk 0.13fF
C1171 ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C1172 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_0/op 0.08fF
C1173 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C1174 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/inv_1/op 0.13fF
C1175 gnd ffipg_3/k 0.61fF
C1176 inv_3/in nand_2/b 0.13fF
C1177 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/op 0.04fF
C1178 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_3/a 0.04fF
C1179 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_0/q 0.20fF
C1180 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_1/a 0.06fF
C1181 ffipg_2/k ffipg_2/ffi_1/q 0.46fF
C1182 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# 0.04fF
C1183 nor_4/b nor_4/a 0.42fF
C1184 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C1185 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C1186 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a 0.00fF
C1187 gnd ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C1188 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_1/b 0.13fF
C1189 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C1190 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C1191 ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C1192 sumffo_0/xor_0/inv_0/op gnd 0.32fF
C1193 ffipg_3/ffi_0/nand_0/w_0_0# ffipg_3/ffi_0/inv_0/op 0.06fF
C1194 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C1195 gnd sumffo_0/ffo_0/nand_0/b 0.58fF
C1196 sumffo_3/xor_0/inv_1/op gnd 0.35fF
C1197 ffipg_1/ffi_0/nand_2/w_0_0# clk 0.06fF
C1198 inv_7/in inv_7/w_0_6# 0.10fF
C1199 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1200 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/q 0.06fF
C1201 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C1202 gnd ffipg_3/ffi_1/inv_1/op 1.85fF
C1203 gnd inv_7/w_0_6# 0.15fF
C1204 y3in gnd 0.22fF
C1205 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C1206 gnd ffipg_0/ffi_0/nand_3/b 0.74fF
C1207 clk sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1208 sumffo_1/sbar z2o 0.32fF
C1209 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_1/b 0.04fF
C1210 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_0/inv_1/op 0.75fF
C1211 sumffo_0/xor_0/w_n3_4# ffi_0/q 0.06fF
C1212 sumffo_3/xor_0/w_n3_4# ffipg_3/k 0.06fF
C1213 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C1214 ffo_0/nand_6/a gnd 0.33fF
C1215 sumffo_3/xor_0/inv_1/w_0_6# gnd 0.06fF
C1216 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a 0.13fF
C1217 gnd cla_2/n 0.60fF
C1218 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k 0.06fF
C1219 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C1220 nor_0/w_0_0# nor_0/a 0.06fF
C1221 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/inv_1/op 0.13fF
C1222 sumffo_0/ffo_0/nand_7/w_0_0# gnd 0.10fF
C1223 ffi_0/nand_1/b ffi_0/nand_7/a 0.13fF
C1224 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C1225 sumffo_2/xor_0/inv_1/op ffi_0/q 0.04fF
C1226 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C1227 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_3/b 0.04fF
C1228 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C1229 gnd ffipg_3/ffi_0/nand_1/b 0.57fF
C1230 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a 0.00fF
C1231 ffipg_3/ffi_1/nand_3/w_0_0# gnd 0.11fF
C1232 nor_4/b gnd 0.25fF
C1233 ffo_0/nand_1/a ffo_0/nand_1/w_0_0# 0.06fF
C1234 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/d 0.06fF
C1235 cla_1/inv_0/in cla_2/p0 0.02fF
C1236 sumffo_1/xor_0/a_38_n43# ffi_0/q 0.01fF
C1237 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/k 0.45fF
C1238 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C1239 y2in ffipg_1/ffi_0/inv_0/op 0.04fF
C1240 ffo_0/nand_3/a ffo_0/nand_3/w_0_0# 0.06fF
C1241 cla_0/l cla_1/n 0.13fF
C1242 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C1243 sumffo_1/ffo_0/inv_0/w_0_6# sumffo_1/ffo_0/inv_0/op 0.03fF
C1244 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b 0.13fF
C1245 ffi_0/nand_6/w_0_0# ffi_0/nand_6/a 0.06fF
C1246 ffipg_2/ffi_1/inv_1/w_0_6# gnd 0.06fF
C1247 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a 0.13fF
C1248 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_1/op 0.06fF
C1249 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C1250 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_1/op 0.52fF
C1251 cla_0/l cla_0/n 0.19fF
C1252 clk ffipg_1/ffi_0/nand_1/a 0.13fF
C1253 ffipg_1/ffi_0/q ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C1254 sumffo_2/ffo_0/nand_0/b clk 0.04fF
C1255 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C1256 cla_0/l cla_2/p0 0.44fF
C1257 inv_3/w_0_6# cla_0/n 0.14fF
C1258 gnd ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C1259 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C1260 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C1261 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C1262 ffo_0/nand_0/b gnd 0.58fF
C1263 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C1264 cla_1/nor_0/w_0_0# gnd 0.31fF
C1265 clk ffi_0/nand_1/a 0.13fF
C1266 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar 0.32fF
C1267 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a 0.31fF
C1268 sumffo_1/xor_0/w_n3_4# ffi_0/q 0.00fF
C1269 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/b 0.31fF
C1270 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_0/q 0.12fF
C1271 ffipg_3/ffi_1/nand_0/w_0_0# ffipg_3/ffi_1/inv_0/op 0.06fF
C1272 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C1273 ffo_0/nand_0/w_0_0# gnd 0.10fF
C1274 sumffo_3/ffo_0/inv_1/w_0_6# gnd 0.06fF
C1275 sumffo_3/ffo_0/nand_6/w_0_0# gnd 0.10fF
C1276 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1277 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1278 cla_1/nand_0/a_13_n26# gnd 0.01fF
C1279 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_1/q 0.06fF
C1280 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_1/b 0.04fF
C1281 ffipg_0/ffi_0/q ffipg_0/ffi_1/q 0.73fF
C1282 gnd sumffo_3/ffo_0/nand_3/b 0.74fF
C1283 gnd ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C1284 ffipg_2/ffi_1/nand_4/w_0_0# gnd 0.10fF
C1285 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/ffi_0/q 0.23fF
C1286 gnd ffo_0/d 0.45fF
C1287 gnd sumffo_3/sbar 0.62fF
C1288 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/ffo_0/nand_6/a 0.06fF
C1289 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C1290 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# 0.04fF
C1291 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C1292 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_4/w_0_0# 0.04fF
C1293 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_1/a 0.06fF
C1294 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/a 0.31fF
C1295 ffipg_0/ffi_1/nand_2/w_0_0# x1in 0.06fF
C1296 sumffo_1/ffo_0/inv_0/w_0_6# sumffo_1/ffo_0/d 0.06fF
C1297 gnd sumffo_0/xor_0/a_10_10# 0.93fF
C1298 cla_2/nor_1/w_0_0# cla_2/g1 0.02fF
C1299 nor_3/b gnd 0.33fF
C1300 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/w_0_0# 0.06fF
C1301 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C1302 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C1303 cla_1/l cla_1/nor_0/w_0_0# 0.05fF
C1304 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C1305 clk ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C1306 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C1307 cla_0/l ffipg_2/k 0.10fF
C1308 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_3/b 0.04fF
C1309 gnd sumffo_2/xor_0/w_n3_4# 0.12fF
C1310 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_3/b 0.31fF
C1311 inv_7/in inv_7/op 0.04fF
C1312 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C1313 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_1/w_0_6# 0.03fF
C1314 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/k 0.45fF
C1315 ffipg_2/ffi_1/nand_0/w_0_0# gnd 0.10fF
C1316 ffipg_1/ffi_1/nand_1/w_0_0# gnd 0.10fF
C1317 ffipg_0/ffi_0/qbar gnd 0.67fF
C1318 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_0/op 0.08fF
C1319 gnd ffo_0/nand_2/w_0_0# 0.10fF
C1320 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/a 0.00fF
C1321 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C1322 sumffo_0/ffo_0/inv_1/w_0_6# sumffo_0/ffo_0/nand_0/b 0.03fF
C1323 inv_7/op gnd 0.27fF
C1324 gnd x2in 0.22fF
C1325 gnd ffipg_0/ffi_0/inv_1/op 1.85fF
C1326 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C1327 ffi_0/nand_7/a ffi_0/nand_5/w_0_0# 0.04fF
C1328 ffipg_1/ffi_0/nand_3/w_0_0# ffipg_1/ffi_0/nand_1/b 0.04fF
C1329 cla_0/l ffipg_1/ffi_0/q 0.13fF
C1330 ffipg_3/ffi_0/inv_1/op y4in 0.01fF
C1331 ffipg_1/ffi_1/inv_0/op ffipg_1/ffi_1/inv_0/w_0_6# 0.03fF
C1332 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a 0.31fF
C1333 inv_8/w_0_6# inv_7/op 0.06fF
C1334 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1335 nor_2/w_0_0# inv_4/in 0.11fF
C1336 gnd ffo_0/nand_3/b 0.74fF
C1337 nor_1/b cla_0/n 0.36fF
C1338 ffi_0/nand_7/w_0_0# ffi_0/q 0.04fF
C1339 gnd ffipg_0/ffi_0/nand_4/w_0_0# 0.10fF
C1340 ffipg_3/ffi_1/inv_0/op x4in 0.04fF
C1341 clk ffipg_2/ffi_0/nand_1/a 0.13fF
C1342 clk ffipg_1/ffi_0/inv_1/op 0.07fF
C1343 cla_1/n gnd 0.51fF
C1344 ffipg_3/ffi_0/q ffipg_3/ffi_1/q 0.73fF
C1345 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1346 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C1347 gnd cla_0/n 0.84fF
C1348 gnd ffi_0/nand_1/w_0_0# 0.10fF
C1349 ffipg_2/pggen_0/nor_0/w_0_0# gnd 0.11fF
C1350 ffipg_2/ffi_1/nand_6/a gnd 0.37fF
C1351 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# 0.04fF
C1352 ffipg_0/ffi_0/nand_2/w_0_0# gnd 0.10fF
C1353 cla_2/p0 gnd 1.06fF
C1354 clk ffipg_3/ffi_1/inv_0/op 0.32fF
C1355 clk ffipg_2/ffi_0/nand_3/a 0.13fF
C1356 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_5/w_0_0# 0.06fF
C1357 ffi_0/nand_3/w_0_0# gnd 0.11fF
C1358 gnd ffipg_0/ffi_1/nand_6/a 0.37fF
C1359 ffi_0/nand_1/b gnd 0.57fF
C1360 ffipg_2/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C1361 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/b 0.31fF
C1362 ffipg_0/ffi_0/inv_0/op gnd 0.27fF
C1363 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C1364 ffipg_2/ffi_1/nand_7/w_0_0# ffipg_2/ffi_1/qbar 0.06fF
C1365 cla_2/p1 ffipg_3/ffi_0/q 0.03fF
C1366 clk ffipg_1/ffi_1/nand_1/a 0.13fF
C1367 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C1368 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C1369 gnd sumffo_2/ffo_0/inv_0/w_0_6# 0.07fF
C1370 z1o sumffo_0/sbar 0.32fF
C1371 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op 0.13fF
C1372 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# 0.04fF
C1373 gnd z4o 0.80fF
C1374 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_3/b 0.00fF
C1375 sumffo_2/ffo_0/nand_4/w_0_0# gnd 0.10fF
C1376 gnd ffipg_3/ffi_0/nand_3/b 0.74fF
C1377 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C1378 sumffo_1/xor_0/a_10_10# ffi_0/q 0.04fF
C1379 gnd cinin 0.22fF
C1380 ffipg_2/ffi_0/nand_1/w_0_0# gnd 0.10fF
C1381 ffipg_0/ffi_0/inv_1/w_0_6# gnd 0.06fF
C1382 clk ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C1383 sumffo_1/ffo_0/nand_7/w_0_0# gnd 0.10fF
C1384 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C1385 ffi_0/inv_1/op ffi_0/inv_1/w_0_6# 0.04fF
C1386 clk ffi_0/inv_0/op 0.32fF
C1387 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C1388 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_0/op 0.06fF
C1389 z3o sumffo_2/ffo_0/nand_7/w_0_0# 0.04fF
C1390 ffipg_3/ffi_0/inv_0/op y4in 0.04fF
C1391 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C1392 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1393 ffipg_0/ffi_1/inv_0/w_0_6# x1in 0.06fF
C1394 ffo_0/nand_1/w_0_0# gnd 0.10fF
C1395 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/sbar 0.06fF
C1396 gnd sumffo_0/ffo_0/nand_1/b 0.57fF
C1397 cla_1/l cla_0/n 0.01fF
C1398 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C1399 clk y1in 0.68fF
C1400 sumffo_1/ffo_0/nand_7/a gnd 0.33fF
C1401 ffipg_3/k ffipg_3/ffi_1/q 0.46fF
C1402 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a 0.00fF
C1403 ffipg_0/ffi_0/q nor_0/a 0.03fF
C1404 ffo_0/nand_3/a ffo_0/nand_0/b 0.13fF
C1405 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/qbar 0.06fF
C1406 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C1407 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C1408 cla_1/l cla_2/p0 0.02fF
C1409 cla_0/l cla_2/l 0.37fF
C1410 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C1411 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a 0.31fF
C1412 ffipg_3/ffi_1/inv_0/w_0_6# x4in 0.06fF
C1413 sumffo_0/xor_0/w_n3_4# sumffo_0/ffo_0/d 0.02fF
C1414 gnd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C1415 ffipg_1/ffi_0/nand_0/w_0_0# gnd 0.10fF
C1416 ffipg_1/ffi_0/q ffipg_1/k 0.07fF
C1417 ffo_0/inv_0/op ffo_0/nand_0/b 0.32fF
C1418 clk ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C1419 ffipg_2/k gnd 0.58fF
C1420 ffipg_0/ffi_0/nand_1/a gnd 0.44fF
C1421 z3o sumffo_2/sbar 0.32fF
C1422 cla_0/inv_0/w_0_6# gnd 0.06fF
C1423 gnd ffi_0/nand_2/w_0_0# 0.10fF
C1424 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/ffi_1/q 0.06fF
C1425 clk ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1426 clk ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C1427 clk sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1428 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1429 ffo_0/inv_0/op ffo_0/nand_0/w_0_0# 0.06fF
C1430 sumffo_2/ffo_0/nand_5/w_0_0# gnd 0.10fF
C1431 cla_2/p1 ffipg_3/k 0.05fF
C1432 gnd ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C1433 cla_1/p0 ffipg_1/ffi_1/q 0.22fF
C1434 cla_1/inv_0/w_0_6# cla_0/n 0.25fF
C1435 ffipg_1/ffi_0/q gnd 3.00fF
C1436 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C1437 ffi_0/nand_3/b gnd 0.74fF
C1438 ffipg_0/ffi_0/nand_6/w_0_0# gnd 0.10fF
C1439 inv_5/in nor_3/b 0.04fF
C1440 ffo_0/inv_0/op ffo_0/d 0.04fF
C1441 cla_0/l cla_0/inv_0/op 0.35fF
C1442 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1443 cla_1/n cla_1/nand_0/w_0_0# 0.04fF
C1444 cla_0/inv_0/in cla_1/p0 0.02fF
C1445 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_1/b 0.04fF
C1446 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a 0.00fF
C1447 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_3/b 0.33fF
C1448 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q 0.22fF
C1449 x3in ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C1450 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/w_0_0# 0.06fF
C1451 sumffo_2/xor_0/inv_1/w_0_6# gnd 0.06fF
C1452 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/q 0.06fF
C1453 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_1/b 0.31fF
C1454 gnd ffipg_1/ffi_1/inv_1/op 1.85fF
C1455 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/w_0_0# 0.06fF
C1456 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C1457 gnd ffipg_3/ffi_1/nand_1/b 0.57fF
C1458 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_6/a 0.04fF
C1459 ffo_0/nand_3/a ffo_0/nand_2/w_0_0# 0.04fF
C1460 sumffo_2/ffo_0/nand_1/b clk 0.45fF
C1461 sumffo_3/xor_0/a_38_n43# ffi_0/q 0.01fF
C1462 cla_0/l cla_0/g0 0.14fF
C1463 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/qbar 0.04fF
C1464 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_5/w_0_0# 0.06fF
C1465 nor_0/b ffi_0/nand_6/w_0_0# 0.04fF
C1466 gnd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C1467 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b 0.13fF
C1468 ffi_0/nand_5/w_0_0# gnd 0.10fF
C1469 ffipg_0/ffi_0/nand_7/w_0_0# gnd 0.10fF
C1470 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C1471 clk ffi_0/inv_1/op 0.93fF
C1472 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C1473 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q 0.32fF
C1474 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# 0.16fF
C1475 nand_2/b cla_0/n 0.00fF
C1476 gnd ffi_0/nand_0/w_0_0# 0.10fF
C1477 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C1478 clk ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C1479 clk ffipg_2/ffi_0/inv_0/op 0.32fF
C1480 gnd ffipg_2/ffi_0/nand_0/a_13_n26# 0.01fF
C1481 ffipg_2/k sumffo_2/xor_0/inv_0/op 0.20fF
C1482 inv_3/in nor_2/b 0.04fF
C1483 nor_2/b inv_4/in 0.16fF
C1484 gnd cla_2/inv_0/op 0.27fF
C1485 inv_5/in cla_0/n 0.13fF
C1486 ffipg_0/ffi_1/nand_2/w_0_0# ffipg_0/ffi_1/nand_3/a 0.04fF
C1487 z3o gnd 0.80fF
C1488 sumffo_0/ffo_0/nand_5/w_0_0# gnd 0.10fF
C1489 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C1490 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C1491 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/a 0.31fF
C1492 nor_4/a inv_8/in 0.04fF
C1493 ffo_0/nand_5/w_0_0# clk 0.06fF
C1494 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C1495 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C1496 clk sumffo_0/ffo_0/nand_3/b 0.33fF
C1497 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/w_0_0# 0.06fF
C1498 gnd ffipg_2/ffi_1/nand_1/w_0_0# 0.10fF
C1499 ffipg_0/pggen_0/xor_0/a_10_10# gnd 0.93fF
C1500 ffi_0/nand_4/w_0_0# ffi_0/inv_1/op 0.06fF
C1501 ffipg_0/ffi_0/nand_3/a gnd 0.33fF
C1502 inv_4/op inv_4/in 0.04fF
C1503 cla_1/p0 nor_0/a 0.24fF
C1504 cla_2/l gnd 0.57fF
C1505 x3in ffipg_2/ffi_1/inv_0/op 0.04fF
C1506 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# 0.04fF
C1507 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C1508 inv_9/in nor_4/w_0_0# 0.11fF
C1509 gnd sumffo_1/ffo_0/inv_0/op 0.27fF
C1510 cla_2/inv_0/w_0_6# gnd 0.06fF
C1511 ffipg_3/ffi_1/nand_3/b gnd 0.74fF
C1512 y4in ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C1513 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# 0.04fF
C1514 ffipg_2/k inv_1/op 0.09fF
C1515 ffipg_0/ffi_0/nand_5/w_0_0# gnd 0.10fF
C1516 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# 0.16fF
C1517 ffo_0/nand_6/a couto 0.31fF
C1518 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a 0.00fF
C1519 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C1520 ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1521 ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1522 ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1523 ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1524 ffipg_3/ffi_1/qbar Gnd 0.42fF
C1525 ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1526 ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1527 ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1528 ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1529 ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1530 ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1531 ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1532 ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1533 x4in Gnd 0.51fF
C1534 ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1535 ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1536 ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1537 ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1538 ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1539 ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1540 ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1541 ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1542 ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1543 ffipg_3/ffi_0/qbar Gnd 0.42fF
C1544 ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1545 ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1546 ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1547 ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1548 ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1549 ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1550 ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1551 ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1552 y4in Gnd 0.51fF
C1553 ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1554 ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1555 ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1556 ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C1557 ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1558 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1559 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1560 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1561 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1562 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1563 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1564 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1565 ffipg_3/ffi_0/q Gnd 2.68fF
C1566 ffipg_3/ffi_1/q Gnd 2.93fF
C1567 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1568 ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1569 ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1570 ffi_0/q Gnd 1.94fF
C1571 ffi_0/nand_7/a Gnd 0.30fF
C1572 ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1573 nor_0/b Gnd 1.01fF
C1574 ffi_0/nand_6/a Gnd 0.30fF
C1575 ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1576 ffi_0/inv_1/op Gnd 0.89fF
C1577 ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1578 ffi_0/nand_3/b Gnd 0.43fF
C1579 ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1580 ffi_0/nand_3/a Gnd 0.30fF
C1581 ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1582 clk Gnd 15.13fF
C1583 cinin Gnd 0.51fF
C1584 ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1585 ffi_0/inv_0/op Gnd 0.26fF
C1586 ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1587 ffi_0/nand_1/a Gnd 0.30fF
C1588 ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1589 ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1590 ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1591 ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C1592 ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1593 ffipg_2/ffi_1/qbar Gnd 0.42fF
C1594 ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C1595 ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1596 ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C1597 ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1598 ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C1599 ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1600 ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C1601 ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1602 x3in Gnd 0.51fF
C1603 ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1604 ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C1605 ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1606 ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C1607 ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1608 ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1609 ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1610 ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C1611 ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1612 ffipg_2/ffi_0/qbar Gnd 0.42fF
C1613 ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C1614 ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1615 ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C1616 ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1617 ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C1618 ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1619 ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C1620 ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1621 y3in Gnd 0.51fF
C1622 ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1623 ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C1624 ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1625 ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C1626 ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1627 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1628 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1629 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1630 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1631 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1632 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1633 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1634 ffipg_2/ffi_0/q Gnd 2.68fF
C1635 ffipg_2/ffi_1/q Gnd 2.93fF
C1636 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1637 ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1638 ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1639 ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C1640 ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1641 ffipg_1/ffi_1/qbar Gnd 0.42fF
C1642 ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C1643 ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1644 ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C1645 ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1646 ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C1647 ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1648 ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C1649 ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1650 x2in Gnd 0.51fF
C1651 ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1652 ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C1653 ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1654 ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C1655 ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1656 ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1657 ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1658 ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C1659 ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1660 ffipg_1/ffi_0/qbar Gnd 0.42fF
C1661 ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C1662 ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1663 ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C1664 ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1665 ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C1666 ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1667 ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C1668 ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1669 y2in Gnd 0.43fF
C1670 ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1671 ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C1672 ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1673 ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C1674 ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1675 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1676 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1677 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1678 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1679 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1680 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1681 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1682 ffipg_1/ffi_0/q Gnd 2.68fF
C1683 ffipg_1/ffi_1/q Gnd 2.93fF
C1684 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1685 inv_9/in Gnd 0.23fF
C1686 nor_4/w_0_0# Gnd 1.81fF
C1687 ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1688 ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1689 ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C1690 ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1691 ffipg_0/ffi_1/qbar Gnd 0.42fF
C1692 ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C1693 ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1694 ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C1695 ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1696 ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C1697 ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1698 ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C1699 ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1700 x1in Gnd 0.39fF
C1701 ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1702 ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C1703 ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1704 ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C1705 ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1706 ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1707 ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1708 ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C1709 ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1710 ffipg_0/ffi_0/qbar Gnd 0.42fF
C1711 ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C1712 ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1713 ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C1714 ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1715 ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C1716 ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1717 ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C1718 ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1719 y1in Gnd 0.51fF
C1720 ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1721 ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C1722 ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1723 ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C1724 ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1725 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1726 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1727 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1728 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1729 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1730 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1731 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1732 ffipg_0/ffi_0/q Gnd 2.68fF
C1733 ffipg_0/ffi_1/q Gnd 2.93fF
C1734 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1735 nor_4/a Gnd 0.43fF
C1736 inv_8/in Gnd 0.22fF
C1737 inv_8/w_0_6# Gnd 1.40fF
C1738 inv_7/in Gnd 0.22fF
C1739 inv_7/w_0_6# Gnd 1.40fF
C1740 inv_5/in Gnd 0.22fF
C1741 inv_5/w_0_6# Gnd 1.40fF
C1742 nor_3/b Gnd 1.17fF
C1743 cla_2/n Gnd 0.36fF
C1744 nor_4/b Gnd 0.32fF
C1745 inv_6/in Gnd 0.23fF
C1746 nor_3/w_0_0# Gnd 1.81fF
C1747 cla_1/n Gnd 0.36fF
C1748 inv_4/in Gnd 0.23fF
C1749 nor_2/w_0_0# Gnd 1.81fF
C1750 nor_2/b Gnd 1.11fF
C1751 inv_3/in Gnd 0.22fF
C1752 inv_3/w_0_6# Gnd 1.40fF
C1753 nor_1/b Gnd 0.91fF
C1754 inv_2/in Gnd 0.22fF
C1755 inv_2/w_0_6# Gnd 1.40fF
C1756 inv_1/in Gnd 0.23fF
C1757 nor_1/w_0_0# Gnd 1.81fF
C1758 inv_0/in Gnd 0.23fF
C1759 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1760 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1761 ffo_0/nand_7/a Gnd 0.30fF
C1762 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1763 ffo_0/qbar Gnd 0.42fF
C1764 ffo_0/nand_6/a Gnd 0.30fF
C1765 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1766 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1767 ffo_0/nand_3/b Gnd 0.43fF
C1768 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1769 ffo_0/nand_3/a Gnd 0.30fF
C1770 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1771 ffo_0/nand_0/b Gnd 0.63fF
C1772 ffo_0/d Gnd 0.42fF
C1773 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1774 ffo_0/inv_0/op Gnd 0.26fF
C1775 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1776 ffo_0/nand_1/a Gnd 0.30fF
C1777 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1778 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1779 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1780 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1781 ffipg_3/k Gnd 1.99fF
C1782 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1783 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1784 inv_4/op Gnd 1.37fF
C1785 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1786 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1787 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1788 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1789 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1790 sumffo_3/sbar Gnd 0.43fF
C1791 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1792 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1793 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1794 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1795 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1796 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1797 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1798 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1799 sumffo_3/ffo_0/d Gnd 0.64fF
C1800 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1801 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1802 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1803 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1804 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1805 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1806 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1807 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1808 nand_2/b Gnd 2.00fF
C1809 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1810 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1811 ffipg_1/k Gnd 2.04fF
C1812 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1813 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1814 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1815 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1816 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1817 sumffo_1/sbar Gnd 0.43fF
C1818 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1819 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1820 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1821 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1822 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1823 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1824 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1825 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1826 sumffo_1/ffo_0/d Gnd 0.64fF
C1827 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1828 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1829 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1830 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1831 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1832 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1833 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1834 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1835 ffipg_2/k Gnd 2.01fF
C1836 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1837 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1838 inv_1/op Gnd 1.37fF
C1839 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1840 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1841 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1842 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1843 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1844 sumffo_2/sbar Gnd 0.43fF
C1845 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1846 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1847 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1848 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1849 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1850 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1851 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1852 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1853 sumffo_2/ffo_0/d Gnd 0.64fF
C1854 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1855 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1856 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1857 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1858 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1859 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1860 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1861 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1862 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1863 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1864 ffipg_0/k Gnd 1.89fF
C1865 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1866 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1867 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1868 gnd Gnd 75.41fF
C1869 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1870 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1871 sumffo_0/sbar Gnd 0.43fF
C1872 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1873 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1874 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1875 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1876 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1877 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1878 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1879 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1880 sumffo_0/ffo_0/d Gnd 0.64fF
C1881 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1882 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1883 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1884 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1885 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1886 cla_2/p1 Gnd 1.09fF
C1887 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1888 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1889 cla_2/inv_0/in Gnd 0.27fF
C1890 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1891 cla_2/g1 Gnd 0.59fF
C1892 cla_2/inv_0/op Gnd 0.26fF
C1893 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1894 cla_1/nor_1/w_0_0# Gnd 1.23fF
C1895 cla_1/l Gnd 0.30fF
C1896 cla_1/nor_0/w_0_0# Gnd 1.23fF
C1897 cla_1/inv_0/in Gnd 0.27fF
C1898 cla_1/inv_0/w_0_6# Gnd 0.58fF
C1899 cla_1/inv_0/op Gnd 0.26fF
C1900 cla_1/nand_0/w_0_0# Gnd 0.82fF
C1901 inv_7/op Gnd 0.26fF
C1902 cla_0/nor_1/w_0_0# Gnd 1.23fF
C1903 cla_0/l Gnd 0.29fF
C1904 cla_0/nor_0/w_0_0# Gnd 1.23fF
C1905 cla_0/inv_0/in Gnd 0.27fF
C1906 cla_0/inv_0/w_0_6# Gnd 0.58fF
C1907 cla_0/inv_0/op Gnd 0.26fF
C1908 cla_0/nand_0/w_0_0# Gnd 0.82fF
C1909 cla_2/l Gnd 0.80fF
C1910 inv_0/op Gnd 0.23fF
C1911 nor_0/w_0_0# Gnd 2.63fF
