magic
tech scmos
timestamp 1618605809
<< nwell >>
rect -3 34 31 40
rect -3 4 59 34
rect 25 -2 59 4
<< ntransistor >>
rect 8 -43 10 -31
rect 18 -43 20 -31
rect 36 -43 38 -31
rect 46 -43 48 -31
<< ptransistor >>
rect 8 10 10 34
rect 18 10 20 34
rect 36 4 38 28
rect 46 4 48 28
<< ndiffusion >>
rect 7 -43 8 -31
rect 10 -43 18 -31
rect 20 -43 21 -31
rect 35 -43 36 -31
rect 38 -43 46 -31
rect 48 -43 49 -31
<< pdiffusion >>
rect 7 10 8 34
rect 10 10 12 34
rect 16 10 18 34
rect 20 10 21 34
rect 35 4 36 28
rect 38 4 40 28
rect 44 4 46 28
rect 48 4 49 28
<< ndcontact >>
rect 3 -43 7 -31
rect 21 -43 25 -31
rect 31 -43 35 -31
rect 49 -43 53 -31
<< pdcontact >>
rect 3 10 7 34
rect 12 10 16 34
rect 21 10 25 34
rect 31 4 35 28
rect 40 4 44 28
rect 49 4 53 28
<< polysilicon >>
rect 8 34 10 37
rect 18 34 20 37
rect 36 28 38 31
rect 46 28 48 31
rect 8 1 10 10
rect 18 0 20 10
rect 8 -31 10 -4
rect 18 -31 20 -5
rect 36 -7 38 4
rect 36 -31 38 -11
rect 46 -18 48 4
rect 46 -31 48 -22
rect 8 -46 10 -43
rect 18 -46 20 -43
rect 36 -46 38 -43
rect 46 -46 48 -43
<< polycontact >>
rect 34 -11 38 -7
rect 45 -22 49 -18
<< metal1 >>
rect -18 44 -9 47
rect -12 43 -9 44
rect -12 40 59 43
rect 3 34 6 40
rect 22 34 25 40
rect -53 14 -50 17
rect -45 15 -42 18
rect -18 15 -6 18
rect -19 -1 -18 0
rect -9 -8 -6 15
rect 32 34 52 37
rect 32 28 35 34
rect 49 28 52 34
rect 13 7 16 10
rect 13 4 31 7
rect 41 -3 44 4
rect 41 -6 58 -3
rect -9 -11 34 -8
rect 55 -17 58 -6
rect 20 -22 45 -19
rect 55 -21 59 -17
rect 20 -24 23 -22
rect -15 -27 23 -24
rect 55 -25 58 -21
rect -53 -40 -50 -37
rect -15 -37 -12 -27
rect 26 -28 58 -25
rect 26 -31 29 -28
rect -45 -40 -42 -37
rect -18 -40 -12 -37
rect 25 -34 31 -31
rect -15 -50 -10 -47
rect 3 -47 6 -43
rect 50 -47 53 -43
rect -5 -50 59 -47
rect -15 -53 -12 -50
rect -18 -56 -12 -53
<< m2contact >>
rect -50 13 -45 18
rect -50 -41 -45 -36
<< pm12contact >>
rect 6 -4 11 1
rect 15 -5 20 0
<< metal2 >>
rect -49 7 -46 13
rect -49 4 -12 7
rect -15 1 -12 4
rect -15 -2 6 1
rect 15 -15 18 -5
rect -48 -18 18 -15
rect -48 -36 -45 -18
<< m123contact >>
rect -42 44 -37 49
rect -42 -9 -37 -4
rect -24 -5 -19 0
rect -10 -50 -5 -45
<< metal3 >>
rect -42 -4 -39 44
rect -19 -5 -7 -2
rect -10 -45 -7 -5
use inv  inv_0
timestamp 1618579805
transform 1 0 -42 0 1 14
box 0 -15 24 33
use inv  inv_1
timestamp 1618579805
transform 1 0 -42 0 1 -41
box 0 -15 24 33
<< labels >>
rlabel metal1 28 -49 28 -49 1 gnd!
rlabel metal1 27 42 27 42 5 vdd!
rlabel metal1 59 -21 59 -17 7 op
rlabel metal1 -10 41 -10 41 1 vdd!
rlabel metal1 -11 -49 -11 -49 1 gnd!
rlabel metal1 -53 -40 -53 -37 3 b
rlabel metal1 -53 14 -53 17 3 a
<< end >>
