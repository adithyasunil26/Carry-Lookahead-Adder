* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 vdd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=216 pd=98 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=108 ps=62
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 vdd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 s1 cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op s1 sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op s1 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 s1 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 vdd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 s3 ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op s3 sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op s3 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 s3 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 s2 nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op s2 sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op s2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 s2 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 vdd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 s4 ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op s4 sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op s4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 s4 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 vdd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in vdd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 vdd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in vdd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in vdd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 vdd y2in cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 cla_1/g0 x2in vdd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_1/g0 y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 vdd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in vdd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in vdd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 vdd y3in cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 cla_0/l x3in vdd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_0/l y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 vdd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in vdd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in vdd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 vdd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in vdd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 vdd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in vdd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in vdd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 cla_2/p0 cla_0/l 0.08fF
C1 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C2 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C3 sumffo_3/xor_0/inv_1/op s4 0.52fF
C4 vdd inv_8/w_0_6# 0.15fF
C5 inv_5/in vdd 0.30fF
C6 vdd ffipg_3/k 0.35fF
C7 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C8 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C9 x1in ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C10 ffipg_1/pggen_0/xor_0/w_n3_4# y2in 0.06fF
C11 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C12 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C13 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C14 nor_2/b nor_2/w_0_0# 0.06fF
C15 x2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C16 cla_2/p1 gnd 0.68fF
C17 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C18 cla_0/inv_0/op nand_2/b 0.09fF
C19 vdd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C20 inv_3/w_0_6# gnd 0.02fF
C21 gnd cla_2/p0 0.68fF
C22 gnd cla_0/nand_0/a_13_n26# 0.00fF
C23 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C24 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C25 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C26 ffipg_2/pggen_0/xor_0/inv_0/op vdd 0.15fF
C27 vdd nor_4/a 0.19fF
C28 inv_0/op cla_0/g0 0.32fF
C29 vdd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C30 vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C31 cla_2/p0 cla_1/l 0.02fF
C32 inv_3/w_0_6# cla_1/l 0.06fF
C33 cla_1/nor_0/w_0_0# cla_0/l 0.01fF
C34 nor_2/b inv_3/in 0.04fF
C35 sumffo_1/xor_0/inv_1/op s2 0.52fF
C36 cla_0/l cla_2/inv_0/in 0.16fF
C37 vdd cla_2/inv_0/op 0.17fF
C38 vdd sumffo_2/xor_0/inv_0/op 0.15fF
C39 sumffo_2/xor_0/inv_0/op s3 0.06fF
C40 nor_0/w_0_0# nand_2/b 0.04fF
C41 inv_1/in nor_1/w_0_0# 0.11fF
C42 vdd sumffo_0/xor_0/inv_1/op 0.15fF
C43 cla_2/p1 y4in 0.03fF
C44 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C45 nor_3/w_0_0# nor_4/b 0.03fF
C46 vdd ffipg_2/k 0.35fF
C47 ffipg_2/pggen_0/xor_0/inv_0/op x3in 0.27fF
C48 sumffo_1/xor_0/a_10_10# cin 0.06fF
C49 ffipg_0/pggen_0/xor_0/inv_0/op gnd 0.17fF
C50 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C51 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# 0.16fF
C52 vdd sumffo_2/xor_0/inv_1/op 0.15fF
C53 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C54 inv_1/in cla_0/n 0.02fF
C55 s3 sumffo_2/xor_0/inv_1/op 0.52fF
C56 nor_1/b inv_2/in 0.04fF
C57 gnd cla_2/inv_0/in 0.30fF
C58 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C59 cla_0/g0 nor_0/a 0.57fF
C60 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C61 nand_2/b cla_0/n 0.06fF
C62 inv_0/in vdd 0.07fF
C63 gnd cla_0/g0 0.70fF
C64 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C65 cla_0/l cin 0.33fF
C66 ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C67 cla_2/l inv_5/w_0_6# 0.08fF
C68 vdd cla_0/inv_0/in 0.05fF
C69 inv_6/in nor_3/w_0_0# 0.11fF
C70 x3in ffipg_2/k 0.46fF
C71 y2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C72 gnd x2in 0.31fF
C73 nor_0/a y1in 0.03fF
C74 gnd y1in 1.62fF
C75 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C76 inv_7/op gnd 0.10fF
C77 vdd sumffo_2/xor_0/a_10_10# 0.93fF
C78 nor_1/b vdd 0.25fF
C79 s3 sumffo_2/xor_0/a_10_10# 0.45fF
C80 inv_3/w_0_6# nor_2/b 0.03fF
C81 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C82 vdd ffipg_3/pggen_0/xor_0/inv_0/op 0.15fF
C83 vdd cla_1/inv_0/op 0.17fF
C84 gnd cin 0.74fF
C85 cla_2/p1 ffipg_3/k 0.05fF
C86 vdd cla_2/g1 0.35fF
C87 vdd inv_7/in 0.30fF
C88 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C89 cla_2/p0 ffipg_3/k 0.06fF
C90 gnd nor_4/b 0.10fF
C91 y2in ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C92 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/k 0.45fF
C93 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/w_n3_4# 0.06fF
C94 x2in ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C95 vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C96 vdd sumffo_1/xor_0/inv_1/op 0.15fF
C97 sumffo_3/xor_0/a_10_10# cin 0.04fF
C98 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# y4in 0.23fF
C99 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C100 cla_0/l cla_0/inv_0/w_0_6# 0.00fF
C101 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C102 cla_1/p0 cla_0/nor_1/w_0_0# 0.06fF
C103 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C104 cla_1/p0 ffipg_1/k 0.05fF
C105 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C106 cla_1/inv_0/w_0_6# vdd 0.06fF
C107 gnd inv_6/in 0.24fF
C108 inv_8/in cin 0.13fF
C109 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C110 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C111 cla_0/inv_0/op cla_1/g0 0.35fF
C112 cla_1/p0 vdd 0.43fF
C113 cla_0/l cla_0/nand_0/w_0_0# 0.00fF
C114 vdd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C115 cin sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C116 gnd x4in 0.31fF
C117 vdd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C118 gnd y2in 1.68fF
C119 inv_6/in nor_3/b 0.16fF
C120 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C121 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C122 ffipg_3/pggen_0/xor_0/inv_1/op y4in 0.22fF
C123 cla_2/p0 ffipg_2/k 0.05fF
C124 nand_2/b inv_2/in 0.34fF
C125 vdd cla_1/nand_0/w_0_0# 0.10fF
C126 vdd cla_2/nor_0/w_0_0# 0.31fF
C127 inv_5/w_0_6# cla_0/n 0.06fF
C128 gnd cla_0/nand_0/w_0_0# 0.01fF
C129 nor_0/w_0_0# cinbar 0.06fF
C130 inv_7/op inv_8/w_0_6# 0.06fF
C131 ffipg_1/k nand_2/b 0.15fF
C132 inv_8/w_0_6# cin 0.06fF
C133 y2in ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C134 vdd inv_1/in 0.09fF
C135 gnd cout 0.10fF
C136 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C137 x4in y4in 0.73fF
C138 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C139 s1 gnd 0.14fF
C140 vdd inv_7/w_0_6# 0.15fF
C141 vdd nand_2/b 0.92fF
C142 nor_4/w_0_0# inv_9/in 0.11fF
C143 cla_1/g0 cla_0/n 0.13fF
C144 cla_1/n cla_0/l 0.13fF
C145 cla_2/g1 cla_2/p1 0.00fF
C146 x2in ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C147 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C148 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k 0.52fF
C149 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C150 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C151 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C152 inv_1/op nor_1/w_0_0# 0.03fF
C153 sumffo_2/xor_0/inv_0/op cin 0.06fF
C154 nor_4/a nor_4/b 0.42fF
C155 cla_1/n gnd 0.24fF
C156 nor_3/w_0_0# nor_3/b 0.06fF
C157 cin sumffo_0/xor_0/inv_1/op 0.22fF
C158 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C159 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C160 inv_4/op inv_4/in 0.04fF
C161 sumffo_3/xor_0/inv_1/op inv_4/op 0.06fF
C162 cla_0/inv_0/in cla_0/g0 0.16fF
C163 ffipg_1/pggen_0/nand_0/a_13_n26# vdd 0.01fF
C164 gnd inv_0/op 0.10fF
C165 nand_2/b inv_3/in 0.13fF
C166 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C167 x4in ffipg_3/k 0.46fF
C168 sumffo_3/xor_0/inv_0/op s4 0.06fF
C169 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C170 cla_2/l cla_0/n 0.32fF
C171 nor_0/a cla_0/l 0.16fF
C172 cin sumffo_2/xor_0/inv_1/op 0.04fF
C173 gnd cla_0/l 1.44fF
C174 cla_1/g0 cla_1/inv_0/in 0.16fF
C175 vdd y3in 0.15fF
C176 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C177 cla_2/g1 cla_2/inv_0/in 0.04fF
C178 inv_0/in cin 0.07fF
C179 cla_1/p0 cla_2/p0 0.24fF
C180 cla_0/l cla_1/l 0.08fF
C181 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C182 sumffo_2/xor_0/inv_1/w_0_6# vdd 0.06fF
C183 vdd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C184 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.24fF
C185 inv_2/w_0_6# inv_2/in 0.10fF
C186 sumffo_2/xor_0/a_38_n43# cin 0.01fF
C187 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C188 y2in ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C189 vdd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C190 vdd ffipg_2/pggen_0/nand_0/a_13_n26# 0.01fF
C191 vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C192 vdd cla_2/n 0.28fF
C193 sumffo_1/xor_0/a_38_n43# cin 0.01fF
C194 ffipg_3/pggen_0/nor_0/w_0_0# x4in 0.06fF
C195 gnd nor_0/a 0.23fF
C196 sumffo_2/xor_0/w_n3_4# ffipg_2/k 0.06fF
C197 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C198 x3in y3in 0.73fF
C199 cin sumffo_2/xor_0/a_10_10# 0.04fF
C200 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C201 sumffo_1/xor_0/inv_0/op s2 0.06fF
C202 vdd inv_4/in 0.09fF
C203 sumffo_3/xor_0/inv_1/op vdd 0.15fF
C204 cla_2/nor_0/w_0_0# cla_2/p0 0.06fF
C205 inv_7/op inv_7/in 0.04fF
C206 gnd cla_1/l 0.18fF
C207 ffipg_0/k cinbar 0.06fF
C208 x3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C209 vdd inv_2/w_0_6# 0.15fF
C210 gnd nor_3/b 0.10fF
C211 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C212 vdd inv_5/w_0_6# 0.15fF
C213 cin sumffo_1/xor_0/inv_1/op 0.04fF
C214 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C215 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C216 cla_1/p0 cla_0/g0 0.38fF
C217 inv_3/w_0_6# nand_2/b 0.06fF
C218 nor_2/b cla_1/n 0.39fF
C219 nor_2/w_0_0# inv_4/in 0.11fF
C220 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.21fF
C221 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C222 ffipg_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C223 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C224 gnd y4in 1.66fF
C225 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C226 cla_1/p0 x2in 0.22fF
C227 gnd inv_8/in 0.13fF
C228 cla_0/n nor_1/w_0_0# 0.06fF
C229 x2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C230 vdd cla_1/g0 0.55fF
C231 cla_0/l cla_1/nor_1/w_0_0# 0.02fF
C232 s1 sumffo_0/xor_0/inv_1/op 0.52fF
C233 vdd cinbar 0.16fF
C234 vdd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C235 ffipg_0/pggen_0/xor_0/a_10_10# y1in 0.12fF
C236 cla_0/l ffipg_3/k 0.10fF
C237 x4in ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C238 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C239 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C240 ffipg_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C241 nand_2/b cla_0/g0 0.13fF
C242 nor_2/b gnd 0.10fF
C243 vdd sumffo_0/xor_0/inv_0/op 0.15fF
C244 vdd inv_9/in 0.09fF
C245 cla_2/p0 y3in 0.03fF
C246 vdd sumffo_1/xor_0/inv_0/op 0.15fF
C247 inv_5/in gnd 0.19fF
C248 gnd ffipg_3/k 0.31fF
C249 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C250 vdd inv_1/op 0.26fF
C251 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C252 vdd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C253 vdd cla_2/l 0.38fF
C254 inv_7/op inv_7/w_0_6# 0.03fF
C255 vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C256 inv_5/in nor_3/b 0.04fF
C257 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_1/op 0.08fF
C258 nand_2/b cin 0.04fF
C259 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C260 vdd sumffo_0/xor_0/a_10_10# 0.93fF
C261 sumffo_3/xor_0/a_10_10# ffipg_3/k 0.12fF
C262 cla_0/l ffipg_2/k 0.04fF
C263 cla_1/p0 y2in 0.03fF
C264 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C265 ffipg_2/pggen_0/xor_0/inv_0/op gnd 0.21fF
C266 y2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C267 gnd nor_4/a 0.21fF
C268 inv_0/in inv_0/op 0.04fF
C269 y4in ffipg_3/k 0.07fF
C270 vdd ffipg_0/pggen_0/nand_0/a_13_n26# 0.01fF
C271 sumffo_3/xor_0/inv_1/w_0_6# vdd 0.06fF
C272 gnd cla_2/inv_0/op 0.10fF
C273 sumffo_2/xor_0/inv_0/op gnd 0.17fF
C274 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C275 inv_8/w_0_6# inv_8/in 0.10fF
C276 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C277 cla_1/nand_0/a_13_n26# gnd 0.01fF
C278 cla_0/inv_0/in cla_0/l 0.14fF
C279 cla_0/inv_0/op vdd 0.17fF
C280 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C281 gnd ffipg_2/k 0.29fF
C282 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C283 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C284 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C285 ffipg_3/pggen_0/nor_0/w_0_0# y4in 0.06fF
C286 inv_0/in nor_0/a 0.02fF
C287 cla_1/g0 cla_2/p0 0.36fF
C288 inv_0/in gnd 0.24fF
C289 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C290 vdd nor_4/w_0_0# 0.15fF
C291 cla_1/inv_0/op cla_0/l 0.35fF
C292 inv_8/in nor_4/a 0.04fF
C293 cla_2/g1 cla_0/l 0.26fF
C294 ffipg_0/k x1in 0.46fF
C295 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C296 cla_0/l inv_7/in 0.13fF
C297 vdd cla_0/nor_0/w_0_0# 0.31fF
C298 vdd nor_0/w_0_0# 0.46fF
C299 vdd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C300 gnd cla_0/inv_0/in 0.30fF
C301 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/k 0.21fF
C302 vdd nor_1/w_0_0# 0.17fF
C303 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C304 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# 0.16fF
C305 nor_1/b gnd 0.10fF
C306 nand_2/b cla_0/nand_0/w_0_0# 0.05fF
C307 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C308 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C309 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.21fF
C310 gnd cla_1/inv_0/op 0.10fF
C311 cla_2/g1 gnd 0.30fF
C312 vdd cla_0/n 0.56fF
C313 gnd inv_7/in 0.13fF
C314 sumffo_3/xor_0/inv_1/op cin 0.04fF
C315 cla_2/p1 cla_2/l 0.02fF
C316 vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C317 inv_2/w_0_6# cin 0.06fF
C318 inv_8/w_0_6# nor_4/a 0.03fF
C319 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C320 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C321 cla_2/l cla_2/p0 0.16fF
C322 cla_1/g0 cla_0/g0 0.14fF
C323 vdd x1in 0.97fF
C324 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/k 0.21fF
C325 cla_1/p0 cla_0/l 0.02fF
C326 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C327 vdd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C328 cin s4 0.16fF
C329 inv_6/in cla_2/n 0.02fF
C330 vdd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C331 ffipg_3/pggen_0/xor_0/inv_0/op y4in 0.20fF
C332 cla_2/g1 y4in 0.13fF
C333 cla_1/nand_0/w_0_0# cla_0/l 0.06fF
C334 cla_1/p0 nor_0/a 0.24fF
C335 cla_1/p0 gnd 0.68fF
C336 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C337 cla_2/nand_0/w_0_0# vdd 0.10fF
C338 vdd cla_1/inv_0/in 0.05fF
C339 cla_1/p0 cla_1/l 0.16fF
C340 vdd sumffo_3/xor_0/inv_0/op 0.15fF
C341 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C342 inv_7/w_0_6# cla_0/l 0.06fF
C343 cla_1/nand_0/w_0_0# gnd 0.01fF
C344 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k 0.06fF
C345 ffipg_0/pggen_0/xor_0/inv_1/op x1in 0.06fF
C346 sumffo_0/xor_0/inv_0/op cin 0.20fF
C347 vdd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C348 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C349 inv_4/op vdd 0.26fF
C350 sumffo_1/xor_0/inv_0/op cin 0.06fF
C351 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C352 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k 0.06fF
C353 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C354 vdd ffipg_0/k 0.33fF
C355 nor_4/b inv_9/in 0.16fF
C356 gnd inv_1/in 0.24fF
C357 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C358 gnd nand_2/b 0.94fF
C359 vdd ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C360 vdd inv_2/in 0.30fF
C361 vdd ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C362 cla_1/g0 y2in 0.13fF
C363 ffipg_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C364 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C365 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C366 inv_4/op nor_2/w_0_0# 0.03fF
C367 nand_2/b cla_1/l 0.31fF
C368 cin sumffo_0/xor_0/a_10_10# 0.12fF
C369 nor_3/w_0_0# cla_2/n 0.06fF
C370 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C371 vdd cla_0/nor_1/w_0_0# 0.31fF
C372 inv_3/w_0_6# cla_0/n 0.16fF
C373 vdd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C374 x1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C375 vdd ffipg_1/k 0.36fF
C376 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C377 cla_0/l y3in 0.13fF
C378 sumffo_2/xor_0/w_n3_4# inv_1/op 0.06fF
C379 cla_1/g0 cla_0/nand_0/w_0_0# 0.06fF
C380 cla_2/g1 cla_2/inv_0/op 0.35fF
C381 x3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C382 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C383 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C384 nor_0/w_0_0# cla_0/g0 0.06fF
C385 cla_1/n inv_4/in 0.02fF
C386 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C387 y3in ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C388 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k 0.52fF
C389 gnd y3in 1.68fF
C390 vdd nor_2/w_0_0# 0.17fF
C391 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C392 x4in ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C393 ffipg_0/k sumffo_0/xor_0/w_n3_4# 0.06fF
C394 vdd x3in 0.93fF
C395 inv_2/w_0_6# cla_0/l 0.06fF
C396 nor_0/w_0_0# cin 0.16fF
C397 ffipg_0/pggen_0/xor_0/inv_0/op x1in 0.27fF
C398 cla_2/p0 cla_1/inv_0/in 0.02fF
C399 nor_4/w_0_0# nor_4/b 0.06fF
C400 inv_9/in cout 0.04fF
C401 vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C402 gnd cla_2/n 0.32fF
C403 s1 sumffo_0/xor_0/inv_0/op 0.06fF
C404 vdd inv_3/in 0.30fF
C405 ffipg_2/pggen_0/nor_0/w_0_0# y3in 0.06fF
C406 ffipg_0/pggen_0/nor_0/w_0_0# x1in 0.06fF
C407 nor_3/b cla_2/n 0.41fF
C408 gnd inv_4/in 0.24fF
C409 sumffo_3/xor_0/inv_1/op gnd 0.20fF
C410 vdd ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C411 y1in ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C412 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C413 cla_1/p0 ffipg_2/k 0.06fF
C414 gnd inv_2/w_0_6# 0.02fF
C415 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C416 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C417 x1in y1in 0.73fF
C418 cla_1/g0 cla_0/l 0.47fF
C419 vdd sumffo_0/xor_0/w_n3_4# 0.12fF
C420 gnd inv_5/w_0_6# 0.26fF
C421 s1 sumffo_0/xor_0/a_10_10# 0.45fF
C422 gnd s4 0.14fF
C423 cla_1/p0 cla_0/inv_0/in 0.02fF
C424 inv_5/w_0_6# nor_3/b 0.17fF
C425 cla_0/inv_0/op cla_0/nand_0/w_0_0# 0.06fF
C426 ffipg_3/pggen_0/xor_0/w_n3_4# x4in 0.06fF
C427 gnd cla_1/g0 0.28fF
C428 nor_0/a cinbar 0.32fF
C429 ffipg_0/pggen_0/xor_0/w_n3_4# x1in 0.06fF
C430 vdd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C431 cla_1/inv_0/w_0_6# cla_1/inv_0/op 0.03fF
C432 vdd cla_2/p1 0.31fF
C433 sumffo_3/xor_0/a_10_10# s4 0.45fF
C434 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k 0.06fF
C435 nand_2/b ffipg_2/k 0.06fF
C436 cin s2 0.27fF
C437 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/k 0.01fF
C438 sumffo_1/xor_0/w_n3_4# s2 0.02fF
C439 vdd cla_2/p0 0.43fF
C440 inv_3/w_0_6# vdd 0.15fF
C441 cla_2/l cla_0/l 0.37fF
C442 nor_4/w_0_0# cout 0.03fF
C443 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/k 0.21fF
C444 gnd sumffo_0/xor_0/inv_0/op 0.21fF
C445 gnd inv_9/in 0.24fF
C446 nor_2/b inv_4/in 0.16fF
C447 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C448 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C449 ffipg_0/k y1in 0.07fF
C450 x3in cla_2/p0 0.22fF
C451 ffipg_2/pggen_0/xor_0/inv_0/op y3in 0.20fF
C452 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C453 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C454 ffipg_3/pggen_0/nand_0/w_0_0# y4in 0.06fF
C455 gnd inv_1/op 0.32fF
C456 sumffo_3/xor_0/inv_1/op ffipg_3/k 0.22fF
C457 nor_1/b inv_1/in 0.16fF
C458 cla_2/l gnd 0.24fF
C459 ffipg_0/k cin 0.19fF
C460 ffipg_1/pggen_0/xor_0/inv_1/op x2in 0.06fF
C461 vdd ffipg_0/pggen_0/xor_0/inv_0/op 0.15fF
C462 ffipg_1/k cla_0/g0 0.06fF
C463 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.02fF
C464 cla_1/nor_0/w_0_0# vdd 0.31fF
C465 vdd cla_2/inv_0/in 0.05fF
C466 inv_3/w_0_6# inv_3/in 0.10fF
C467 cla_2/l nor_3/b 0.10fF
C468 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C469 vdd cla_0/g0 0.53fF
C470 inv_7/w_0_6# inv_7/in 0.10fF
C471 inv_5/in inv_5/w_0_6# 0.10fF
C472 cla_0/inv_0/op cla_0/l 0.21fF
C473 cin inv_2/in 0.13fF
C474 y3in ffipg_2/k 0.07fF
C475 ffipg_1/k x2in 0.46fF
C476 ffipg_0/pggen_0/nor_0/w_0_0# vdd 0.11fF
C477 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C478 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/k 0.02fF
C479 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C480 nor_0/w_0_0# inv_0/op 0.10fF
C481 vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C482 vdd x2in 0.93fF
C483 sumffo_2/xor_0/inv_1/w_0_6# ffipg_2/k 0.23fF
C484 ffipg_1/k cin 0.06fF
C485 vdd y1in 0.15fF
C486 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C487 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C488 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C489 inv_7/op vdd 0.17fF
C490 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C491 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C492 vdd cin 0.78fF
C493 cla_0/inv_0/op gnd 0.10fF
C494 vdd sumffo_1/xor_0/w_n3_4# 0.12fF
C495 cin s3 0.28fF
C496 cin sumffo_3/xor_0/a_38_n43# 0.01fF
C497 vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C498 vdd nor_4/b 0.15fF
C499 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C500 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C501 cla_2/inv_0/w_0_6# vdd 0.06fF
C502 cla_0/l cla_0/n 0.12fF
C503 vdd ffipg_3/pggen_0/xor_0/inv_1/op 0.15fF
C504 nor_0/w_0_0# nor_0/a 0.06fF
C505 cla_2/p1 cla_2/p0 0.24fF
C506 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C507 ffipg_0/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C508 vdd ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C509 ffipg_1/pggen_0/xor_0/inv_1/op y2in 0.22fF
C510 vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C511 x3in ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C512 sumffo_2/xor_0/w_n3_4# s3 0.02fF
C513 inv_5/in cla_2/l 0.05fF
C514 cla_2/g1 cla_2/n 0.13fF
C515 vdd inv_6/in 0.09fF
C516 ffipg_0/pggen_0/xor_0/inv_1/op y1in 0.22fF
C517 ffipg_1/k y2in 0.07fF
C518 cla_1/g0 ffipg_2/k 0.06fF
C519 gnd cla_0/n 0.61fF
C520 vdd cla_0/inv_0/w_0_6# 0.06fF
C521 vdd x4in 0.93fF
C522 nor_1/b inv_2/w_0_6# 0.03fF
C523 vdd y2in 0.15fF
C524 nor_4/a inv_9/in 0.02fF
C525 sumffo_1/xor_0/a_10_10# s2 0.45fF
C526 cla_1/l cla_0/n 0.07fF
C527 ffipg_3/pggen_0/xor_0/w_n3_4# y4in 0.06fF
C528 x1in nor_0/a 0.22fF
C529 gnd x1in 0.22fF
C530 cla_2/p1 cla_2/inv_0/in 0.02fF
C531 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C532 inv_0/in cinbar 0.16fF
C533 cin sumffo_0/xor_0/w_n3_4# 0.06fF
C534 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C535 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C536 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C537 cla_1/g0 cla_0/inv_0/in 0.04fF
C538 gnd sumffo_0/xor_0/inv_0/w_0_6# 0.02fF
C539 cla_0/l cla_1/inv_0/in 0.07fF
C540 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C541 vdd cla_0/nand_0/w_0_0# 0.10fF
C542 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C543 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C544 vdd cout 0.15fF
C545 ffipg_0/pggen_0/nand_0/w_0_0# y1in 0.06fF
C546 inv_1/op ffipg_2/k 0.09fF
C547 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C548 gnd s2 0.14fF
C549 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C550 cla_2/nand_0/w_0_0# gnd 0.08fF
C551 gnd cla_1/inv_0/in 0.30fF
C552 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C553 vdd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C554 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C555 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C556 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/k 0.02fF
C557 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C558 ffipg_3/pggen_0/xor_0/a_10_10# y4in 0.12fF
C559 vdd nor_3/w_0_0# 0.14fF
C560 cla_0/l cla_0/nor_1/w_0_0# 0.00fF
C561 inv_4/op gnd 0.32fF
C562 vdd cla_1/n 0.28fF
C563 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C564 ffipg_0/k nor_0/a 0.05fF
C565 nor_4/w_0_0# nor_4/a 0.07fF
C566 vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C567 gnd ffipg_0/k 0.41fF
C568 inv_5/in cla_0/n 0.13fF
C569 cla_0/n ffipg_3/k 0.06fF
C570 vdd sumffo_1/xor_0/a_10_10# 0.93fF
C571 vdd inv_0/op 0.17fF
C572 ffipg_0/pggen_0/xor_0/inv_0/op y1in 0.20fF
C573 cla_1/p0 cla_1/g0 0.07fF
C574 cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C575 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C576 cla_0/g0 y1in 0.13fF
C577 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C578 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C579 gnd inv_2/in 0.17fF
C580 vdd cla_0/l 1.05fF
C581 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.24fF
C582 cla_1/n nor_2/w_0_0# 0.06fF
C583 cla_0/g0 cin 0.08fF
C584 inv_2/w_0_6# nand_2/b 0.03fF
C585 cla_2/p1 x4in 0.22fF
C586 ffipg_0/pggen_0/nor_0/w_0_0# y1in 0.06fF
C587 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C588 vdd ffipg_2/pggen_0/xor_0/inv_1/op 0.15fF
C589 ffipg_1/k nor_0/a 0.06fF
C590 s1 sumffo_0/xor_0/w_n3_4# 0.02fF
C591 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C592 ffipg_1/k gnd 0.39fF
C593 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/k 0.45fF
C594 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C595 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C596 vdd cla_2/nor_1/w_0_0# 0.31fF
C597 gnd cla_2/nand_0/a_13_n26# 0.01fF
C598 vdd nor_0/a 0.35fF
C599 vdd gnd 3.73fF
C600 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C601 inv_7/op cin 0.31fF
C602 inv_0/in nor_0/w_0_0# 0.11fF
C603 gnd s3 0.14fF
C604 y3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C605 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C606 sumffo_3/xor_0/w_n3_4# s4 0.02fF
C607 vdd cla_1/l 0.22fF
C608 cin sumffo_1/xor_0/w_n3_4# 0.00fF
C609 y3in ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C610 cla_1/g0 nand_2/b 0.06fF
C611 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C612 x3in ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C613 vdd nor_3/b 0.23fF
C614 ffipg_2/k cla_0/n 0.06fF
C615 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C616 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C617 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C618 ffipg_1/pggen_0/xor_0/w_n3_4# x2in 0.06fF
C619 sumffo_3/xor_0/a_10_10# vdd 0.93fF
C620 ffipg_0/pggen_0/xor_0/w_n3_4# y1in 0.06fF
C621 vdd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C622 x3in gnd 0.31fF
C623 vdd ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C624 nor_1/b nor_1/w_0_0# 0.06fF
C625 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C626 vdd y4in 0.10fF
C627 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C628 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C629 inv_4/op ffipg_3/k 0.09fF
C630 sumffo_2/xor_0/w_n3_4# cin 0.00fF
C631 vdd inv_8/in 0.30fF
C632 gnd inv_3/in 0.17fF
C633 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C634 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C635 y2in x2in 0.73fF
C636 inv_1/in inv_1/op 0.04fF
C637 vdd sumffo_0/xor_0/inv_1/w_0_6# 0.07fF
C638 ffipg_0/pggen_0/xor_0/inv_1/op gnd 0.20fF
C639 nor_1/b cla_0/n 0.36fF
C640 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C641 inv_7/w_0_6# cla_2/l 0.06fF
C642 cla_1/inv_0/op cla_0/n 0.06fF
C643 inv_6/in nor_4/b 0.04fF
C644 cla_2/p1 cla_0/l 0.30fF
C645 nor_2/b vdd 0.21fF
C646 vdd cla_1/nor_1/w_0_0# 0.31fF
C647 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C648 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C649 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C650 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C651 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C652 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C653 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C654 y4in Gnd 2.72fF
C655 x4in Gnd 2.80fF
C656 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C657 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C658 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C659 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C660 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C661 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C662 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C663 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C664 y3in Gnd 2.72fF
C665 x3in Gnd 2.80fF
C666 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C667 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C668 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C669 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C670 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C671 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C672 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C673 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C674 y2in Gnd 2.72fF
C675 x2in Gnd 2.80fF
C676 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C677 cout Gnd 0.19fF
C678 inv_9/in Gnd 0.23fF
C679 nor_4/w_0_0# Gnd 1.81fF
C680 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C681 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C682 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C683 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C684 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C685 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C686 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C687 y1in Gnd 2.72fF
C688 x1in Gnd 2.80fF
C689 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C690 nor_4/a Gnd 0.59fF
C691 inv_8/in Gnd 0.22fF
C692 inv_8/w_0_6# Gnd 1.40fF
C693 inv_7/in Gnd 0.22fF
C694 inv_7/w_0_6# Gnd 1.40fF
C695 nor_4/b Gnd 0.32fF
C696 nor_3/b Gnd 0.77fF
C697 inv_5/in Gnd 0.22fF
C698 inv_5/w_0_6# Gnd 1.40fF
C699 cla_2/n Gnd 0.36fF
C700 inv_6/in Gnd 0.23fF
C701 nor_3/w_0_0# Gnd 1.81fF
C702 vdd Gnd 8.88fF
C703 cla_1/n Gnd 0.36fF
C704 inv_4/in Gnd 0.23fF
C705 nor_2/w_0_0# Gnd 1.81fF
C706 cla_0/n Gnd 1.34fF
C707 nor_2/b Gnd 0.82fF
C708 inv_3/in Gnd 0.22fF
C709 inv_3/w_0_6# Gnd 1.40fF
C710 cinbar Gnd 1.21fF
C711 nor_0/a Gnd 2.07fF
C712 nor_1/b Gnd 1.05fF
C713 inv_2/in Gnd 0.22fF
C714 inv_2/w_0_6# Gnd 1.40fF
C715 inv_1/in Gnd 0.23fF
C716 nor_1/w_0_0# Gnd 1.81fF
C717 inv_0/in Gnd 0.23fF
C718 s4 Gnd 0.07fF
C719 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C720 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C721 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C722 ffipg_3/k Gnd 2.89fF
C723 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C724 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C725 inv_4/op Gnd 1.37fF
C726 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C727 s2 Gnd 0.07fF
C728 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C729 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C730 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C731 nand_2/b Gnd 2.36fF
C732 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C733 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C734 ffipg_1/k Gnd 2.78fF
C735 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C736 s3 Gnd 0.07fF
C737 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C738 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C739 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C740 ffipg_2/k Gnd 2.89fF
C741 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C742 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C743 inv_1/op Gnd 1.30fF
C744 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C745 s1 Gnd 0.07fF
C746 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C747 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C748 gnd Gnd 23.13fF
C749 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C750 cin Gnd 7.80fF
C751 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C752 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C753 ffipg_0/k Gnd 1.49fF
C754 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C755 cla_2/p1 Gnd 1.09fF
C756 cla_2/nor_1/w_0_0# Gnd 1.23fF
C757 cla_2/nor_0/w_0_0# Gnd 1.23fF
C758 cla_2/inv_0/in Gnd 0.27fF
C759 cla_2/inv_0/w_0_6# Gnd 0.58fF
C760 cla_2/g1 Gnd 0.59fF
C761 cla_2/inv_0/op Gnd 0.26fF
C762 cla_2/nand_0/w_0_0# Gnd 0.82fF
C763 cla_2/p0 Gnd 0.38fF
C764 cla_1/nor_1/w_0_0# Gnd 1.23fF
C765 cla_1/l Gnd 0.30fF
C766 cla_1/nor_0/w_0_0# Gnd 1.23fF
C767 cla_1/inv_0/in Gnd 0.27fF
C768 cla_1/inv_0/w_0_6# Gnd 0.58fF
C769 cla_1/inv_0/op Gnd 0.26fF
C770 cla_1/nand_0/w_0_0# Gnd 0.82fF
C771 inv_7/op Gnd 0.26fF
C772 cla_1/p0 Gnd 2.28fF
C773 cla_0/nor_1/w_0_0# Gnd 1.23fF
C774 cla_0/l Gnd 1.95fF
C775 cla_0/nor_0/w_0_0# Gnd 1.23fF
C776 cla_0/inv_0/in Gnd 0.27fF
C777 cla_0/inv_0/w_0_6# Gnd 0.58fF
C778 cla_1/g0 Gnd 1.49fF
C779 cla_0/inv_0/op Gnd 0.26fF
C780 cla_0/nand_0/w_0_0# Gnd 0.82fF
C781 cla_2/l Gnd 0.25fF
C782 cla_0/g0 Gnd 1.40fF
C783 inv_0/op Gnd 0.23fF
C784 nor_0/w_0_0# Gnd 2.63fF
