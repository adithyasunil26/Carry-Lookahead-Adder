magic
tech scmos
timestamp 1618844298
<< metal1 >>
rect -3 1270 97 1273
rect 102 1270 802 1273
rect 3 1263 666 1266
rect 3 1256 6 1263
rect -3 1252 0 1255
rect 241 1212 533 1215
rect 241 1156 497 1159
rect -3 1153 0 1156
rect -3 1083 0 1086
rect 479 1014 484 1019
rect 494 998 497 1156
rect 530 1148 533 1212
rect 530 1145 549 1148
rect 671 1143 674 1146
rect 897 1137 900 1140
rect 539 1026 542 1036
rect 563 1023 572 1026
rect 970 1001 971 1004
rect 494 995 505 998
rect 563 994 572 997
rect 606 993 618 996
rect 490 989 505 992
rect 566 988 572 991
rect 566 966 569 988
rect 490 963 576 966
rect 611 939 618 942
rect -3 876 0 879
rect 611 874 614 939
rect 481 871 614 874
rect -3 802 0 805
rect 481 738 484 871
rect 479 735 484 738
rect -3 595 0 598
rect -3 521 0 524
rect -3 314 0 317
rect -3 237 0 240
rect -2 30 1 33
rect -2 -8 40 -5
rect 45 -8 569 -5
<< metal2 >>
rect 481 1199 552 1202
rect 481 1019 484 1199
rect 479 1014 484 1019
rect 479 735 484 738
<< m123contact >>
rect 97 1270 102 1275
rect 802 1269 807 1274
rect 666 1261 671 1266
rect 666 1143 671 1148
rect 539 1036 544 1041
rect 537 970 542 975
rect 576 963 581 968
rect 40 -9 45 -4
<< metal3 >>
rect 98 1245 101 1270
rect 667 1148 670 1261
rect 803 1229 806 1269
rect 699 1056 702 1164
rect 757 1072 760 1112
rect 757 1069 832 1072
rect 699 1053 775 1056
rect 407 1043 542 1046
rect 407 1030 410 1043
rect 539 1041 542 1043
rect 772 982 775 1053
rect 829 1034 832 1069
rect 539 966 542 970
rect 539 963 576 966
rect 539 937 542 963
rect 449 934 542 937
rect 41 -4 44 46
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 548 0 1 1105
box -3 -9 349 129
use nor  nor_0
timestamp 1618580541
transform 1 0 505 0 1 1000
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 539 0 1 993
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 572 0 1 999
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1618628987
transform 1 0 621 0 -1 1036
box -3 -9 349 129
<< labels >>
rlabel metal1 -3 314 -3 317 3 y3in
rlabel metal1 -3 1153 -3 1156 3 cinin
rlabel metal1 -3 1083 -3 1086 3 x1in
rlabel metal1 -3 876 -3 879 3 y1in
rlabel metal1 -3 802 -3 805 3 x2in
rlabel metal1 -3 595 -3 598 3 y2in
rlabel metal1 -3 521 -3 524 3 x3in
rlabel metal1 -3 237 -3 240 3 x4in
rlabel metal1 -2 30 -2 33 3 y4in
rlabel metal1 -3 1252 -3 1255 3 clk
rlabel metal1 71 1271 71 1271 5 vdd!
rlabel metal1 19 -7 19 -7 1 gnd!
rlabel metal1 900 1137 900 1140 7 z1o
rlabel metal1 971 1001 971 1004 7 z2o
<< end >>
