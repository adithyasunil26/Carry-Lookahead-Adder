magic
tech scmos
timestamp 1618628828
<< metal1 >>
rect 110 120 135 123
rect -3 94 -2 97
rect 122 91 128 94
rect 122 62 125 91
rect 348 88 349 91
rect 110 59 125 62
rect -3 40 -2 43
rect 126 38 127 41
rect 348 32 349 35
<< m2contact >>
rect 135 54 140 59
rect 107 30 112 35
<< metal2 >>
rect 109 54 135 57
rect 109 35 112 54
use xor  xor_0
timestamp 1618605809
transform 1 0 51 0 1 80
box -53 -56 59 49
use ffo  ffo_0
timestamp 1618618535
transform 1 0 141 0 1 33
box -14 -42 207 91
<< labels >>
rlabel metal1 349 32 349 35 7 q
rlabel metal1 349 88 349 91 7 qbar
rlabel metal1 -3 94 -3 97 3 k
rlabel metal1 -3 40 -3 43 3 c
rlabel metal1 126 38 126 41 1 clk
<< end >>
