`timescale 1ns / 1ps

`include "cla.v"

module clatb;

  reg clk ;
  reg x1  ;
  reg x2  ;
  reg x3  ;
  reg x4  ;
  reg y1  ;
  reg y2  ;
  reg y3  ;
  reg y4  ;
  reg cin ;
  
  wire z1  ;
  wire z2  ;
  wire z3  ;
  wire z4  ;
  wire cout;

  
  cla cla1(
    .x1   (x1  ) ,
    .x2   (x2  ) ,
    .x3   (x3  ) ,
    .x4   (x4  ) ,
    .y1   (y1  ) ,
    .y2   (y2  ) ,
    .y3   (y3  ) ,
    .y4   (y4  ) ,
    .cin  (cin ) ,
    .z1   (z1  ) ,
    .z2   (z2  ) ,
    .z3   (z3  ) ,
    .z4   (z4  ) ,
    .cout (cout)
  );

  reg [4:1] x;
  reg [4:1] y;
  reg [4:1] z;

  initial begin 
    $dumpfile("test.vcd");
    $dumpvars(0,clatb);
    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 0; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 0; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 0; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 0; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 0; y3  = 1; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 0;    
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 0; y2  = 1; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 0; y1  = 1; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 0; cin = 1;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 0;
    #5 clk = 0; #5 clk = 1; x4  = 1; x3  = 1; x2  = 1; x1  = 1; y4  = 1; y3  = 1; y2  = 1; y1  = 1; cin = 1;      

  end 

  always@(posedge clk)
  begin
    x={x4,x3,x2,x1};
    y={y4,y3,y2,y1};
    z={z4,z3,z2,z1};
  end

  initial 
		// $monitor("clk=%b x1=%b x2=%b x3=%b x4=%b y1=%b y2=%b y3=%b y4=%b cin=%b z1=%b z2=%b z3=%b z4=%b cout=%b",clk,x1,x2,x3,x4,y1,y2,y3,y4,cin,z1,z2,z3,z4,cout);
    $monitor("clk=%d x=%d y=%d cin=%d z=%d cout=%d",clk,x,y,cin,z,cout);
endmodule
