* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 vdd a_13_n18# a_10_10# w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1005 op a_13_n18# a_10_n43# Gnd nfet w=12 l=2
+  ad=192 pd=56 as=96 ps=40
M1006 gnd inv_1/op a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1007 a_10_10# inv_1/op op w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1008 a_10_n43# a gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_38_n43# inv_0/op op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_10_10# a vdd w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 op inv_0/op a_10_10# w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b inv_1/op 0.09fF
C1 inv_0/w_0_6# a 0.06fF
C2 gnd b 0.05fF
C3 inv_0/op vdd 0.15fF
C4 op w_n3_4# 0.02fF
C5 a vdd 0.11fF
C6 vdd inv_1/in 0.02fF
C7 b a_13_n18# 0.09fF
C8 vdd inv_1/op 0.15fF
C9 gnd vdd 0.25fF
C10 op inv_0/op 0.06fF
C11 op inv_1/op 0.50fF
C12 vdd a_10_10# 0.93fF
C13 op gnd 0.10fF
C14 inv_1/in inv_1/w_0_6# 0.06fF
C15 inv_1/op inv_1/w_0_6# 0.03fF
C16 vdd b 0.10fF
C17 op a_10_10# 0.45fF
C18 inv_0/w_0_6# vdd 0.09fF
C19 inv_0/op w_n3_4# 0.06fF
C20 a w_n3_4# 0.06fF
C21 w_n3_4# inv_1/op 0.06fF
C22 b inv_1/w_0_6# 0.17fF
C23 a inv_0/op 0.27fF
C24 w_n3_4# a_13_n18# 0.06fF
C25 inv_0/op inv_1/op 0.08fF
C26 inv_0/op gnd 0.17fF
C27 w_n3_4# a_10_10# 0.16fF
C28 a inv_1/op 0.06fF
C29 vdd inv_1/w_0_6# 0.06fF
C30 a gnd 0.22fF
C31 inv_1/in inv_1/op 0.04fF
C32 gnd inv_1/in 0.05fF
C33 inv_0/op a_13_n18# 0.06fF
C34 gnd inv_1/op 0.20fF
C35 a a_13_n18# 0.02fF
C36 inv_1/op a_13_n18# 0.12fF
C37 inv_0/op b 0.07fF
C38 w_n3_4# vdd 0.12fF
C39 a b 0.00fF
C40 inv_0/w_0_6# inv_0/op 0.03fF
C41 a_10_10# a_13_n18# 0.06fF
C42 inv_1/in b 0.00fF
C43 b Gnd 0.61fF **FLOATING
C44 op Gnd 0.03fF
C45 a_10_10# Gnd 0.01fF
C46 a_13_n18# Gnd 0.27fF
C47 w_n3_4# Gnd 1.14fF
C48 gnd Gnd 0.72fF
C49 inv_1/op Gnd 0.49fF
C50 vdd Gnd 0.59fF
C51 inv_1/in Gnd 0.14fF
C52 inv_1/w_0_6# Gnd 0.58fF
C53 inv_0/op Gnd 0.51fF
C54 a Gnd 1.25fF
C55 inv_0/w_0_6# Gnd 0.58fF
