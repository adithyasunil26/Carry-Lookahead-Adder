magic
tech scmos
timestamp 1618833724
<< metal1 >>
rect 0 1270 97 1273
rect 102 1270 525 1273
rect 3 1263 632 1266
rect 3 1256 6 1263
rect 241 1212 423 1215
rect 420 1165 423 1212
rect 420 1162 514 1165
rect 639 1160 643 1163
rect 866 1154 869 1157
rect 490 989 498 992
rect 490 963 491 966
rect 518 732 519 735
rect 490 708 519 711
rect 487 674 490 682
rect 518 680 519 683
rect 487 671 519 674
rect 501 643 504 671
rect 515 451 519 454
rect 490 427 519 430
rect 487 393 490 401
rect 518 399 519 402
rect 487 390 519 393
rect 501 374 504 390
rect 490 143 519 146
rect 487 109 490 117
rect 517 115 519 118
rect 487 106 519 109
rect 22 -13 73 -10
rect 78 -13 233 -10
<< m2contact >>
rect 498 987 503 992
rect 491 961 496 966
rect 513 732 518 737
rect 513 680 518 685
rect 500 638 505 643
rect 513 399 518 404
rect 500 369 505 374
rect 514 167 519 172
rect 512 115 517 120
<< metal2 >>
rect 478 1216 518 1219
rect 478 1019 481 1216
rect 481 653 484 706
rect 492 683 495 961
rect 500 735 503 987
rect 500 732 513 735
rect 492 680 513 683
rect 481 650 518 653
rect 481 383 484 425
rect 501 402 504 638
rect 515 451 518 650
rect 501 399 513 402
rect 481 380 519 383
rect 501 118 504 369
rect 516 172 519 380
rect 501 115 512 118
<< m123contact >>
rect 97 1270 102 1275
rect 525 1270 530 1275
rect 632 1261 637 1266
rect 634 1160 639 1165
rect 563 773 568 778
rect 600 651 605 656
rect 563 492 568 497
rect 600 370 605 375
rect 563 208 568 213
rect 600 86 605 91
rect 73 -14 78 -9
<< metal3 >>
rect 98 1245 101 1270
rect 526 1251 529 1270
rect 634 1165 637 1261
rect 408 780 566 783
rect 408 749 411 780
rect 563 778 566 780
rect 449 653 600 656
rect 408 499 566 502
rect 408 468 411 499
rect 563 497 566 499
rect 449 372 600 375
rect 408 216 566 219
rect 408 184 411 216
rect 563 213 566 216
rect 449 88 600 91
rect 74 -9 77 58
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 517 0 1 1122
box -3 -9 349 129
use cla  cla_0
timestamp 1618627066
transform 1 0 528 0 1 683
box -9 -46 112 95
use cla  cla_1
timestamp 1618627066
transform 1 0 528 0 1 402
box -9 -46 112 95
use cla  cla_2
timestamp 1618627066
transform 1 0 528 0 1 118
box -9 -46 112 95
<< labels >>
rlabel metal1 869 1154 869 1157 7 z1o
<< end >>
