* SPICE3 file created from ffipgarrcla.ext - technology: scmos

.option scale=0.09u

M1000 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=7410 ps=4464
M1001 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=14820 pd=8198 as=96 ps=40
M1002 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1005 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1006 cla_0/l cla_0/p0 cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1007 cla_0/nor_0/a_13_6# cla_0/p1 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 gnd cla_0/p0 cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1009 cla_0/l cla_0/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1011 cla_0/nor_1/a_13_6# cla_0/p1 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1013 cla_0/inv_0/in cla_0/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1015 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1016 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1018 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1019 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1021 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1023 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1025 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1027 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1029 vdd ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1030 cla_0/g0 ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 cla_0/g0 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1032 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1033 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1034 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1035 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1036 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1037 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1038 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1039 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1040 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 cla_0/p0 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd ffipgarr_0/ffipg_0/ffi_1/q cla_0/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_0/p0 ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1049 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1050 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1052 ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 ffipgarr_0/ffipg_0/ffi_0/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# ffipgarr_0/y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1057 vdd sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1058 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/y1in vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 ffipgarr_0/ffipg_0/ffi_0/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1060 ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1061 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1062 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1064 ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1065 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1066 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1069 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1070 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1072 ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1073 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1074 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1076 ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1077 vdd ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1078 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/y1in vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 ffipgarr_0/ffipg_0/ffi_0/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1083 ffipgarr_0/ffipg_0/ffi_0/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1084 ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1086 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1088 ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1089 vdd sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1090 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 ffipgarr_0/ffipg_0/ffi_1/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# ffipgarr_0/x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 vdd sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1094 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/x1in vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 ffipgarr_0/ffipg_0/ffi_1/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1096 ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1097 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1098 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1101 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1102 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1105 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1106 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1108 ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1109 vdd ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1110 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1112 ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1113 vdd ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1114 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/x1in vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 ffipgarr_0/ffipg_0/ffi_1/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 ffipgarr_0/ffipg_0/ffi_1/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 vdd ffipgarr_0/ffipg_1/ffi_0/q cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1122 cla_1/g0 ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1124 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1127 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1128 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1129 ffipgarr_0/k2 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1130 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1131 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1132 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/k2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 cla_0/p1 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1137 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 gnd ffipgarr_0/ffipg_1/ffi_1/q cla_0/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1139 cla_0/p1 ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1141 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1142 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1145 vdd sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1146 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 ffipgarr_0/ffipg_1/ffi_0/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# ffipgarr_0/y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1149 vdd sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1150 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/y2in vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 ffipgarr_0/ffipg_1/ffi_0/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1157 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1158 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1161 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1162 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1163 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1164 ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1165 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1166 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1168 ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1169 vdd ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1170 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1172 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/y2in vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipgarr_0/ffipg_1/ffi_0/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1175 ffipgarr_0/ffipg_1/ffi_0/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1176 ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1177 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1178 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1181 vdd sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1182 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 ffipgarr_0/ffipg_1/ffi_1/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1184 ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# ffipgarr_0/x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1185 vdd sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1186 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/x2in vdd ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipgarr_0/ffipg_1/ffi_1/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1188 ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1189 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1190 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1192 ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1193 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1194 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1197 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1198 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1201 vdd ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1202 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1204 ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1205 vdd ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1206 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1208 ffipgarr_0/ffipg_1/ffi_1/inv_0/op ffipgarr_0/x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1209 ffipgarr_0/ffipg_1/ffi_1/inv_0/op ffipgarr_0/x2in vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1210 ffipgarr_0/ffipg_1/ffi_1/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1211 ffipgarr_0/ffipg_1/ffi_1/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1212 ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1213 vdd ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1214 cla_2/g0 ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 cla_2/g0 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1216 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1217 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1221 ffipgarr_0/k3 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1222 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1223 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/k3 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1224 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/k3 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipgarr_0/k3 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1229 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 gnd ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1231 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1233 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1234 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1236 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1237 vdd sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1238 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 ffipgarr_0/ffipg_2/ffi_0/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1240 ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# ffipgarr_0/y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1241 vdd sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1242 ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/y3in vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 ffipgarr_0/ffipg_2/ffi_0/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1245 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1246 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1248 ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1249 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1250 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1252 ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1253 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1254 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1256 ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1257 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1258 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1260 ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1261 vdd ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1262 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1264 ffipgarr_0/ffipg_2/ffi_0/inv_0/op ffipgarr_0/y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1265 ffipgarr_0/ffipg_2/ffi_0/inv_0/op ffipgarr_0/y3in vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1266 ffipgarr_0/ffipg_2/ffi_0/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1267 ffipgarr_0/ffipg_2/ffi_0/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1268 ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1269 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1270 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1272 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1273 vdd sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1274 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 ffipgarr_0/ffipg_2/ffi_1/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1276 ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# ffipgarr_0/x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1277 vdd sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1278 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/x3in vdd ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 ffipgarr_0/ffipg_2/ffi_1/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1280 ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1281 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1282 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1284 ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1285 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1286 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1288 ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1289 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1290 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1291 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1293 vdd ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1294 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1297 vdd ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1298 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1301 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/x3in vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1302 ffipgarr_0/ffipg_2/ffi_1/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1303 ffipgarr_0/ffipg_2/ffi_1/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1304 ffipgarr_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1305 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1306 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/a vdd ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1308 ffipgarr_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1309 vdd sumffo_0/clk ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1310 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/inv_0/op vdd ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 ffipgarr_0/ffi_0/nand_1/a sumffo_0/clk ffipgarr_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 ffipgarr_0/ffi_0/nand_2/a_13_n26# ffipgarr_0/cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1313 vdd sumffo_0/clk ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1314 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/cinin vdd ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 ffipgarr_0/ffi_0/nand_3/a sumffo_0/clk ffipgarr_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1316 ffipgarr_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1317 vdd ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1318 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/a vdd ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1320 ffipgarr_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1321 vdd ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1322 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_3/b vdd ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 ffipgarr_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1325 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1326 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/inv_1/op vdd ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1328 ffipgarr_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1329 vdd sumffo_0/c ffipgarr_0/cinbar ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1330 ffipgarr_0/cinbar ffipgarr_0/ffi_0/nand_6/a vdd ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 ffipgarr_0/cinbar sumffo_0/c ffipgarr_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipgarr_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 vdd ffipgarr_0/cinbar sumffo_0/c ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 sumffo_0/c ffipgarr_0/ffi_0/nand_7/a vdd ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 sumffo_0/c ffipgarr_0/cinbar ffipgarr_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1337 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/cinin vdd ffipgarr_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1338 ffipgarr_0/ffi_0/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1339 ffipgarr_0/ffi_0/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1341 vdd ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1342 cla_2/g1 ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1344 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1345 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1346 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1347 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1348 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1349 ffipgarr_0/k4 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1350 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1351 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/k4 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1352 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1353 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/k4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 ffipgarr_0/k4 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1356 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1357 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 gnd ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1359 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1360 ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1361 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1362 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 vdd sumffo_0/clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 ffipgarr_0/ffipg_3/ffi_0/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# ffipgarr_0/y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1369 vdd sumffo_0/clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1370 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/y4in vdd ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1371 ffipgarr_0/ffipg_3/ffi_0/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1373 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1374 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1376 ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1377 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1378 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1380 ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1381 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1382 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1384 ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1385 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1386 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 vdd ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1393 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/y4in vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1394 ffipgarr_0/ffipg_3/ffi_0/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1395 ffipgarr_0/ffipg_3/ffi_0/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 vdd sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipgarr_0/ffipg_3/ffi_1/nand_1/a sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# ffipgarr_0/x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 vdd sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/x4in vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipgarr_0/ffipg_3/ffi_1/nand_3/a sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1417 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1418 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1421 vdd ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1422 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1425 vdd ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1426 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1427 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1428 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1429 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/x4in vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1430 ffipgarr_0/ffipg_3/ffi_1/inv_1/op sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1431 ffipgarr_0/ffipg_3/ffi_1/inv_1/op sumffo_0/clk vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1433 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1434 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1436 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1437 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1438 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1439 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1441 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1443 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1445 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1447 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1448 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a vdd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1450 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1451 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1452 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op vdd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1455 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1456 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1458 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1459 vdd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1460 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a vdd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1463 vdd sumffo_0/clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1464 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b vdd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 sumffo_0/ffo_0/nand_6/a sumffo_0/clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1466 sumffo_0/ffo_0/nand_5/a_13_n26# sumffo_0/clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1467 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1468 sumffo_0/ffo_0/nand_7/a sumffo_0/clk vdd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1470 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 vdd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a vdd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 vdd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 z1o sumffo_0/ffo_0/nand_7/a vdd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1480 sumffo_0/ffo_0/nand_0/b sumffo_0/clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1481 sumffo_0/ffo_0/nand_0/b sumffo_0/clk vdd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 sumffo_0/xor_0/inv_0/op sumffo_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1483 sumffo_0/xor_0/inv_0/op sumffo_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1484 sumffo_0/xor_0/inv_1/op sumffo_0/c gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1485 sumffo_0/xor_0/inv_1/op sumffo_0/c vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 vdd sumffo_0/c sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1487 sumffo_0/ffo_0/d sumffo_0/c sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1488 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1489 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1490 sumffo_0/xor_0/a_10_n43# sumffo_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1491 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 sumffo_0/xor_0/a_10_10# sumffo_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C1 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C2 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C3 ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C4 ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C5 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C6 ffipgarr_0/ffipg_2/ffi_0/q gnd 2.62fF
C7 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C8 sumffo_0/c ffipgarr_0/ffi_0/nand_7/w_0_0# 0.04fF
C9 ffipgarr_0/ffi_0/nand_7/w_0_0# vdd 0.10fF
C10 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C11 gnd ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.15fF
C12 ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd 0.34fF
C13 vdd sumffo_0/ffo_0/nand_6/a 0.30fF
C14 cla_2/p1 cla_2/inv_0/in 0.02fF
C15 ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd 0.39fF
C16 ffipgarr_0/ffi_0/inv_1/w_0_6# ffipgarr_0/ffi_0/inv_1/op 0.04fF
C17 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C18 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.04fF
C19 sumffo_0/k sumffo_0/xor_0/w_n3_4# 0.06fF
C20 ffipgarr_0/ffi_0/nand_3/b vdd 0.39fF
C21 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.04fF
C22 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.32fF
C23 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# vdd 0.10fF
C24 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.04fF
C25 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C26 ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd 0.03fF
C27 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# sumffo_0/clk 0.06fF
C28 gnd sumffo_0/ffo_0/nand_6/a 0.03fF
C29 ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd 0.35fF
C30 ffipgarr_0/k3 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C31 ffipgarr_0/cinbar ffipgarr_0/ffi_0/nand_6/w_0_0# 0.04fF
C32 ffipgarr_0/ffi_0/inv_0/op vdd 0.17fF
C33 ffipgarr_0/ffi_0/nand_3/b gnd 0.35fF
C34 cla_0/p0 sumffo_0/k 0.05fF
C35 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C36 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# vdd 0.10fF
C37 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C38 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# vdd 0.93fF
C39 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# vdd 0.10fF
C40 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/q 0.00fF
C41 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C42 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C43 cla_0/g0 vdd 0.40fF
C44 cla_0/p0 cla_0/l 0.16fF
C45 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/q 0.00fF
C46 cla_2/g0 cla_2/inv_0/in 0.16fF
C47 vdd sumffo_0/ffo_0/nand_0/w_0_0# 0.10fF
C48 ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd 0.30fF
C49 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C50 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# cla_0/p1 0.24fF
C51 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C52 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_0/q 0.12fF
C53 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.75fF
C54 ffipgarr_0/ffi_0/inv_0/op gnd 0.10fF
C55 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# vdd 0.10fF
C56 ffipgarr_0/ffi_0/inv_1/op sumffo_0/clk 0.10fF
C57 sumffo_0/c vdd 0.38fF
C58 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_0/q 0.73fF
C59 cla_1/inv_0/in cla_1/inv_0/op 0.04fF
C60 ffipgarr_0/ffipg_1/ffi_1/qbar vdd 0.33fF
C61 gnd cla_0/g0 0.03fF
C62 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.04fF
C63 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C64 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# vdd 0.10fF
C65 ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd 0.03fF
C66 ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd 0.30fF
C67 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.13fF
C68 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.04fF
C69 ffipgarr_0/ffipg_3/ffi_0/nand_1/b vdd 0.31fF
C70 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C71 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C72 cla_0/p1 cla_0/g0 0.30fF
C73 ffipgarr_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffi_0/inv_0/op 0.06fF
C74 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C75 sumffo_0/c gnd 0.63fF
C76 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/b 0.31fF
C77 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C78 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/a 0.00fF
C79 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# vdd 0.06fF
C80 ffipgarr_0/ffipg_1/ffi_1/qbar gnd 0.34fF
C81 gnd vdd 3.65fF
C82 ffipgarr_0/x4in ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C83 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.00fF
C84 sumffo_0/ffo_0/nand_3/b vdd 0.39fF
C85 ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd 1.63fF
C86 ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd 0.14fF
C87 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.06fF
C88 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C89 cla_1/g0 cla_0/nand_0/w_0_0# 0.06fF
C90 gnd ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.26fF
C91 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C92 cla_0/p1 vdd 0.37fF
C93 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.13fF
C94 ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd 0.17fF
C95 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# vdd 0.06fF
C96 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# ffipgarr_0/y2in 0.06fF
C97 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C98 ffipgarr_0/ffi_0/nand_0/w_0_0# vdd 0.10fF
C99 ffipgarr_0/ffipg_2/ffi_0/nand_1/b vdd 0.31fF
C100 ffipgarr_0/y1in vdd 0.04fF
C101 sumffo_0/ffo_0/nand_3/b gnd 0.35fF
C102 ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd 0.22fF
C103 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C104 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/q 0.31fF
C105 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.13fF
C106 cla_1/g0 cla_2/p0 0.30fF
C107 gnd ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C108 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/k3 0.52fF
C109 cla_1/inv_0/w_0_6# vdd 0.06fF
C110 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C111 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.00fF
C112 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.03fF
C113 gnd cla_0/p1 1.03fF
C114 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C115 ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd 0.10fF
C116 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.13fF
C117 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C118 sumffo_0/ffo_0/inv_0/w_0_6# sumffo_0/ffo_0/d 0.06fF
C119 gnd ffipgarr_0/ffi_0/nand_0/a_13_n26# 0.01fF
C120 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C121 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/q 0.00fF
C122 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/qbar 0.00fF
C123 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C124 ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd 0.17fF
C125 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a 0.00fF
C126 ffipgarr_0/ffi_0/nand_0/w_0_0# gnd 0.00fF
C127 ffipgarr_0/ffi_0/nand_3/a vdd 0.30fF
C128 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C129 ffipgarr_0/ffipg_2/ffi_0/nand_1/b gnd 0.26fF
C130 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/y2in 0.01fF
C131 gnd ffipgarr_0/y1in 0.19fF
C132 ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C133 ffipgarr_0/ffi_0/nand_1/a vdd 0.30fF
C134 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.45fF
C135 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.32fF
C136 ffipgarr_0/y4in sumffo_0/clk 0.64fF
C137 ffipgarr_0/ffipg_3/ffi_1/nand_1/b vdd 0.31fF
C138 ffipgarr_0/y3in vdd 0.04fF
C139 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# 0.04fF
C140 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.06fF
C141 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C142 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# vdd 0.10fF
C143 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C144 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C145 ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd 0.10fF
C146 ffipgarr_0/ffi_0/nand_3/a gnd 0.03fF
C147 ffipgarr_0/ffi_0/nand_1/a gnd 0.14fF
C148 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/k4 0.01fF
C149 ffipgarr_0/ffi_0/inv_0/w_0_6# ffipgarr_0/ffi_0/inv_0/op 0.03fF
C150 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/a 0.06fF
C151 ffipgarr_0/cinin ffipgarr_0/ffi_0/nand_2/w_0_0# 0.06fF
C152 sumffo_0/clk sumffo_0/ffo_0/nand_1/b 0.45fF
C153 ffipgarr_0/ffipg_3/ffi_1/nand_1/b gnd 0.26fF
C154 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# vdd 0.10fF
C155 ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd 0.17fF
C156 ffipgarr_0/y3in gnd 0.19fF
C157 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/y3in 0.01fF
C158 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C159 cla_0/p0 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C160 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.06fF
C161 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.04fF
C162 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.04fF
C163 sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d 0.06fF
C164 ffipgarr_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffi_0/nand_1/a 0.04fF
C165 ffipgarr_0/x3in ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C166 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C167 ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd 1.63fF
C168 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# vdd 0.10fF
C169 sumffo_0/clk ffipgarr_0/x1in 0.70fF
C170 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# gnd 0.00fF
C171 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C172 cla_0/inv_0/in cla_0/g0 0.16fF
C173 gnd ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.10fF
C174 ffipgarr_0/ffipg_0/ffi_0/qbar vdd 0.33fF
C175 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C176 sumffo_0/sbar vdd 0.28fF
C177 ffipgarr_0/ffipg_3/ffi_0/qbar vdd 0.33fF
C178 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_1/q 0.73fF
C179 ffipgarr_0/ffi_0/inv_0/w_0_6# vdd 0.06fF
C180 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.13fF
C181 ffipgarr_0/ffipg_0/ffi_1/q cla_0/p0 0.22fF
C182 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C183 cla_2/inv_0/op cla_2/nand_0/w_0_0# 0.06fF
C184 cla_2/g0 cla_1/g0 0.10fF
C185 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C186 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/k4 0.02fF
C187 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.04fF
C188 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.00fF
C189 cla_2/g1 vdd 0.35fF
C190 ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd 0.22fF
C191 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.00fF
C192 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C193 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q 0.22fF
C194 ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd 0.34fF
C195 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a 0.13fF
C196 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.75fF
C197 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C198 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C199 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# ffipgarr_0/x1in 0.06fF
C200 gnd ffipgarr_0/ffipg_0/ffi_0/qbar 0.34fF
C201 cla_0/inv_0/in vdd 0.05fF
C202 gnd sumffo_0/sbar 0.34fF
C203 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_0/op 0.32fF
C204 ffipgarr_0/ffipg_3/ffi_0/qbar gnd 0.34fF
C205 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C206 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.06fF
C207 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# vdd 0.10fF
C208 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# sumffo_0/clk 0.06fF
C209 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op vdd 0.15fF
C210 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C211 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# vdd 0.10fF
C212 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.04fF
C213 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# vdd 0.10fF
C214 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/w_0_0# 0.06fF
C215 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C216 ffipgarr_0/y4in ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.01fF
C217 gnd cla_2/g1 0.23fF
C218 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C219 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_6/w_0_0# 0.06fF
C220 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# vdd 0.10fF
C221 gnd ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.03fF
C222 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C223 gnd cla_0/inv_0/in 0.35fF
C224 sumffo_0/ffo_0/nand_7/a vdd 0.30fF
C225 sumffo_0/xor_0/w_n3_4# sumffo_0/ffo_0/d 0.02fF
C226 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# vdd 0.10fF
C227 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.07fF
C228 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C229 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.04fF
C230 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# gnd 0.00fF
C231 cla_2/inv_0/w_0_6# vdd 0.06fF
C232 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op gnd 0.17fF
C233 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/k4 0.46fF
C234 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# sumffo_0/clk 0.06fF
C235 cla_0/p1 cla_0/inv_0/in 0.02fF
C236 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C237 ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd 0.34fF
C238 cla_1/p0 vdd 0.06fF
C239 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# vdd 0.06fF
C240 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.31fF
C241 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.06fF
C242 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.04fF
C243 sumffo_0/ffo_0/nand_7/a gnd 0.03fF
C244 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# vdd 0.10fF
C245 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.07fF
C246 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C247 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.20fF
C248 ffipgarr_0/ffipg_1/ffi_0/qbar vdd 0.33fF
C249 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# vdd 0.10fF
C250 ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd 0.30fF
C251 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# vdd 0.10fF
C252 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_0/q 0.23fF
C253 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.00fF
C254 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# vdd 0.93fF
C255 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.06fF
C256 gnd ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.03fF
C257 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.13fF
C258 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# vdd 0.93fF
C259 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/k4 0.07fF
C260 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.31fF
C261 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/k2 0.02fF
C262 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C263 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.04fF
C264 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/nand_7/a 0.04fF
C265 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# vdd 0.10fF
C266 ffipgarr_0/ffipg_1/ffi_0/qbar gnd 0.34fF
C267 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/q 0.00fF
C268 z1o sumffo_0/ffo_0/nand_6/a 0.31fF
C269 cla_1/p0 cla_0/p1 0.03fF
C270 cla_0/p0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C271 ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd 0.14fF
C272 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C273 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.04fF
C274 ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd 0.39fF
C275 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C276 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/k3 0.01fF
C277 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# vdd 0.10fF
C278 ffipgarr_0/k2 vdd 0.13fF
C279 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op vdd 0.15fF
C280 cla_2/n vdd 0.28fF
C281 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op vdd 0.15fF
C282 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q 0.32fF
C283 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/q 0.04fF
C284 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C285 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C286 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# vdd 0.10fF
C287 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.13fF
C288 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# 0.04fF
C289 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# ffipgarr_0/y1in 0.06fF
C290 cla_2/g0 cla_1/n 0.13fF
C291 ffipgarr_0/k4 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C292 ffipgarr_0/y2in vdd 0.04fF
C293 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.04fF
C294 gnd ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.35fF
C295 ffipgarr_0/ffipg_2/ffi_1/nand_1/b vdd 0.31fF
C296 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C297 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C298 ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 0.22fF
C299 ffipgarr_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C300 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# 0.06fF
C301 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k 0.52fF
C302 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# vdd 0.10fF
C303 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/q 0.00fF
C304 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.00fF
C305 ffipgarr_0/k2 gnd 0.14fF
C306 ffipgarr_0/ffipg_0/ffi_0/q cla_0/p0 0.03fF
C307 gnd cla_2/n 0.03fF
C308 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.75fF
C309 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op gnd 0.20fF
C310 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op gnd 0.20fF
C311 ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd 0.34fF
C312 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# gnd 0.00fF
C313 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/q 0.00fF
C314 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.32fF
C315 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q 0.32fF
C316 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.00fF
C317 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/qbar 0.00fF
C318 ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd 0.39fF
C319 ffipgarr_0/y2in gnd 0.19fF
C320 ffipgarr_0/k2 cla_0/p1 0.05fF
C321 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C322 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# ffipgarr_0/y3in 0.06fF
C323 ffipgarr_0/ffipg_2/ffi_1/nand_1/b gnd 0.26fF
C324 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C325 cla_1/n cla_1/nand_0/w_0_0# 0.04fF
C326 cla_0/nor_1/w_0_0# cla_0/g0 0.06fF
C327 cla_1/g0 cla_0/n 0.13fF
C328 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C329 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# cla_2/p0 0.05fF
C330 z1o vdd 0.28fF
C331 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C332 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.13fF
C333 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C334 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.13fF
C335 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C336 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C337 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.00fF
C338 ffipgarr_0/ffipg_3/ffi_0/q cla_2/p1 0.03fF
C339 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C340 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C341 ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd 0.03fF
C342 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/qbar 0.04fF
C343 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C344 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C345 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C346 ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd 0.30fF
C347 sumffo_0/ffo_0/nand_1/w_0_0# vdd 0.10fF
C348 ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd 0.34fF
C349 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# vdd 0.10fF
C350 ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd 0.35fF
C351 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.45fF
C352 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C353 sumffo_0/ffo_0/nand_7/a sumffo_0/sbar 0.31fF
C354 ffipgarr_0/cinin sumffo_0/clk 0.70fF
C355 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.33fF
C356 ffipgarr_0/ffipg_1/ffi_0/q vdd 0.38fF
C357 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C358 cla_0/nor_1/w_0_0# vdd 0.31fF
C359 gnd z1o 0.52fF
C360 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C361 ffipgarr_0/ffi_0/nand_3/w_0_0# vdd 0.11fF
C362 ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd 0.03fF
C363 sumffo_0/xor_0/inv_1/op sumffo_0/c 0.22fF
C364 ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd 0.03fF
C365 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.32fF
C366 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# 0.04fF
C367 sumffo_0/xor_0/inv_1/op vdd 0.15fF
C368 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C369 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.32fF
C370 gnd cla_0/nor_1/w_0_0# 0.01fF
C371 ffipgarr_0/ffipg_3/ffi_0/nand_3/a sumffo_0/clk 0.13fF
C372 ffipgarr_0/ffipg_1/ffi_0/q gnd 2.62fF
C373 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# vdd 0.06fF
C374 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# vdd 0.06fF
C375 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.04fF
C376 ffipgarr_0/k4 cla_2/p1 0.05fF
C377 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.04fF
C378 ffipgarr_0/ffipg_1/ffi_0/q cla_0/p1 0.03fF
C379 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.06fF
C380 cla_0/p1 cla_0/nor_1/w_0_0# 0.06fF
C381 vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C382 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C383 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C384 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# vdd 0.06fF
C385 cla_1/inv_0/in vdd 0.05fF
C386 gnd cla_1/nor_1/a_13_6# 0.01fF
C387 sumffo_0/xor_0/inv_1/op gnd 0.20fF
C388 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C389 ffipgarr_0/x4in sumffo_0/clk 0.70fF
C390 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.03fF
C391 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# cla_2/g1 0.04fF
C392 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.06fF
C393 sumffo_0/ffo_0/nand_4/w_0_0# vdd 0.10fF
C394 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.06fF
C395 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# 0.06fF
C396 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# vdd 0.10fF
C397 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.03fF
C398 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/qbar 0.31fF
C399 cla_1/nor_1/w_0_0# cla_1/g0 0.06fF
C400 sumffo_0/ffo_0/nand_3/a vdd 0.30fF
C401 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar 0.32fF
C402 ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd 0.34fF
C403 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C404 gnd cla_1/inv_0/in 0.35fF
C405 cla_2/p0 cla_2/p1 0.24fF
C406 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C407 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# ffipgarr_0/y1in 0.06fF
C408 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C409 ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd 1.63fF
C410 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C411 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C412 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C413 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.04fF
C414 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.45fF
C415 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.04fF
C416 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.16fF
C417 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.04fF
C418 ffipgarr_0/ffi_0/nand_2/w_0_0# vdd 0.10fF
C419 sumffo_0/ffo_0/nand_3/a gnd 0.03fF
C420 ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd 0.03fF
C421 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.13fF
C422 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a 0.31fF
C423 cla_2/n cla_2/g1 0.13fF
C424 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.06fF
C425 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.04fF
C426 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C427 ffipgarr_0/x2in ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.01fF
C428 sumffo_0/ffo_0/nand_0/b vdd 0.15fF
C429 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# vdd 0.11fF
C430 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.33fF
C431 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b 0.32fF
C432 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C433 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.13fF
C434 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# vdd 0.10fF
C435 gnd ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.22fF
C436 cla_1/inv_0/in cla_1/inv_0/w_0_6# 0.06fF
C437 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.07fF
C438 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C439 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.06fF
C440 cla_2/g0 cla_2/p0 0.14fF
C441 ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd 0.34fF
C442 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.13fF
C443 z1o sumffo_0/sbar 0.32fF
C444 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# vdd 0.11fF
C445 ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 0.22fF
C446 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.13fF
C447 cla_2/inv_0/in vdd 0.05fF
C448 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_0/qbar 0.06fF
C449 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.13fF
C450 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C451 cla_0/inv_0/w_0_6# vdd 0.06fF
C452 gnd sumffo_0/ffo_0/nand_0/b 0.38fF
C453 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.04fF
C454 ffipgarr_0/x2in ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C455 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/y1in 0.01fF
C456 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.31fF
C457 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/qbar 0.04fF
C458 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.04fF
C459 ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd 0.03fF
C460 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.06fF
C461 ffipgarr_0/ffi_0/nand_1/w_0_0# vdd 0.10fF
C462 cla_2/p0 cla_2/l 0.16fF
C463 vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C464 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.00fF
C465 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C466 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d 0.04fF
C467 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# vdd 0.10fF
C468 gnd cla_2/inv_0/in 0.35fF
C469 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C470 cla_1/l vdd 0.20fF
C471 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.06fF
C472 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.13fF
C473 ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd 0.30fF
C474 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C475 sumffo_0/c sumffo_0/k 0.15fF
C476 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# sumffo_0/clk 0.06fF
C477 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.07fF
C478 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_2/w_0_0# 0.04fF
C479 cla_2/g0 cla_2/p1 0.30fF
C480 ffipgarr_0/ffi_0/nand_1/b vdd 0.31fF
C481 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.04fF
C482 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C483 vdd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C484 sumffo_0/k vdd 0.25fF
C485 cla_0/nor_1/w_0_0# cla_0/inv_0/in 0.05fF
C486 cla_1/g0 cla_0/inv_0/op 0.35fF
C487 sumffo_0/ffo_0/nand_7/a z1o 0.00fF
C488 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.06fF
C489 cla_0/l vdd 0.20fF
C490 gnd cla_1/l 0.18fF
C491 ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd 0.17fF
C492 ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd 0.14fF
C493 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.31fF
C494 ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd 0.34fF
C495 gnd ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C496 ffipgarr_0/ffi_0/nand_7/w_0_0# ffipgarr_0/cinbar 0.06fF
C497 ffipgarr_0/ffi_0/nand_1/b gnd 0.26fF
C498 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.06fF
C499 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C500 gnd sumffo_0/k 0.35fF
C501 cla_2/p1 cla_2/l 0.02fF
C502 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# vdd 0.11fF
C503 gnd cla_0/l 0.18fF
C504 ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd 0.10fF
C505 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C506 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/cinin 0.01fF
C507 ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd 0.03fF
C508 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# vdd 0.10fF
C509 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C510 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C511 cla_0/l cla_0/p1 0.02fF
C512 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# vdd 0.10fF
C513 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/clk 0.06fF
C514 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.13fF
C515 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op vdd 0.15fF
C516 sumffo_0/ffo_0/inv_0/w_0_6# sumffo_0/ffo_0/inv_0/op 0.03fF
C517 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_1/a 0.06fF
C518 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q 0.32fF
C519 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C520 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C521 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/x1in 0.01fF
C522 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C523 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# vdd 0.06fF
C524 gnd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.00fF
C525 cla_2/g0 cla_1/nand_0/w_0_0# 0.06fF
C526 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.17fF
C527 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/a 0.31fF
C528 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.04fF
C529 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.13fF
C530 sumffo_0/clk sumffo_0/ffo_0/nand_6/a 0.13fF
C531 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# cla_1/g0 0.04fF
C532 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C533 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.04fF
C534 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.31fF
C535 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C536 ffipgarr_0/ffipg_0/ffi_0/nand_1/b vdd 0.31fF
C537 ffipgarr_0/ffi_0/inv_1/w_0_6# vdd 0.06fF
C538 cla_1/nor_0/w_0_0# vdd 0.31fF
C539 sumffo_0/c ffipgarr_0/cinbar 0.32fF
C540 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.04fF
C541 ffipgarr_0/x2in vdd 0.04fF
C542 ffipgarr_0/cinbar vdd 0.28fF
C543 ffipgarr_0/y3in ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.04fF
C544 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# vdd 0.11fF
C545 ffipgarr_0/k2 ffipgarr_0/ffipg_1/ffi_0/q 0.07fF
C546 cla_1/g0 cla_0/g0 0.10fF
C547 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# vdd 0.10fF
C548 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# 0.04fF
C549 gnd ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.26fF
C550 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q 0.22fF
C551 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# 0.06fF
C552 sumffo_0/clk ffipgarr_0/ffi_0/inv_0/op 0.32fF
C553 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.04fF
C554 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/qbar 0.31fF
C555 ffipgarr_0/x3in vdd 0.04fF
C556 ffipgarr_0/x2in gnd 0.19fF
C557 ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd 0.34fF
C558 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.06fF
C559 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.04fF
C560 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C561 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C562 cla_2/g1 cla_2/inv_0/in 0.04fF
C563 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C564 ffipgarr_0/cinbar gnd 0.34fF
C565 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.04fF
C566 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.06fF
C567 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.04fF
C568 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C569 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.13fF
C570 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/d 0.06fF
C571 ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd 0.17fF
C572 sumffo_0/c sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C573 cla_1/g0 vdd 0.47fF
C574 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.31fF
C575 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# ffipgarr_0/x3in 0.06fF
C576 sumffo_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C577 ffipgarr_0/x3in gnd 0.19fF
C578 ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd 0.03fF
C579 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C580 cla_2/g0 cla_1/inv_0/op 0.35fF
C581 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.06fF
C582 ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd 0.39fF
C583 sumffo_0/clk vdd 7.21fF
C584 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# vdd 0.10fF
C585 sumffo_0/xor_0/a_10_10# sumffo_0/ffo_0/d 0.45fF
C586 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.13fF
C587 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C588 ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd 0.10fF
C589 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# vdd 0.11fF
C590 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/x3in 0.04fF
C591 ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd 0.34fF
C592 gnd cla_1/g0 0.26fF
C593 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C594 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# ffipgarr_0/y3in 0.06fF
C595 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C596 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.31fF
C597 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# vdd 0.06fF
C598 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.04fF
C599 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# vdd 0.10fF
C600 ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd 0.35fF
C601 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.04fF
C602 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C603 cla_0/p1 cla_1/g0 0.14fF
C604 cla_0/p0 cla_0/nor_0/w_0_0# 0.06fF
C605 sumffo_0/clk gnd 7.22fF
C606 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C607 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.00fF
C608 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.13fF
C609 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C610 sumffo_0/ffo_0/nand_3/b sumffo_0/clk 0.33fF
C611 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# ffipgarr_0/k3 0.21fF
C612 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# vdd 0.06fF
C613 ffipgarr_0/ffipg_0/ffi_1/q vdd 1.31fF
C614 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# vdd 0.10fF
C615 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.07fF
C616 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.33fF
C617 ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd 0.03fF
C618 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C619 sumffo_0/c ffipgarr_0/ffi_0/nand_7/a 0.00fF
C620 ffipgarr_0/ffipg_2/ffi_1/inv_0/op sumffo_0/clk 0.32fF
C621 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C622 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# sumffo_0/k 0.02fF
C623 ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd 0.39fF
C624 ffipgarr_0/ffi_0/nand_7/a vdd 0.30fF
C625 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C626 cla_1/p0 cla_1/l 0.16fF
C627 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# vdd 0.10fF
C628 sumffo_0/ffo_0/inv_1/w_0_6# vdd 0.06fF
C629 cla_2/nand_0/w_0_0# vdd 0.10fF
C630 ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd 0.30fF
C631 sumffo_0/clk ffipgarr_0/y1in 0.70fF
C632 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# vdd 0.10fF
C633 ffipgarr_0/ffi_0/nand_0/w_0_0# sumffo_0/clk 0.06fF
C634 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# vdd 0.06fF
C635 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/x1in 0.04fF
C636 gnd ffipgarr_0/ffipg_0/ffi_1/q 0.93fF
C637 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C638 ffipgarr_0/y4in ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C639 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_4/w_0_0# 0.06fF
C640 ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd 0.30fF
C641 sumffo_0/ffo_0/nand_7/w_0_0# vdd 0.10fF
C642 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C643 gnd ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.35fF
C644 ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd 0.30fF
C645 ffipgarr_0/ffi_0/nand_7/a gnd 0.03fF
C646 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C647 ffipgarr_0/k3 cla_2/p0 0.05fF
C648 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# vdd 0.10fF
C649 ffipgarr_0/ffipg_3/ffi_0/inv_0/op sumffo_0/clk 0.32fF
C650 ffipgarr_0/ffi_0/nand_3/a sumffo_0/clk 0.13fF
C651 ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd 0.03fF
C652 cla_2/nor_1/w_0_0# cla_2/g0 0.06fF
C653 ffipgarr_0/ffi_0/nand_1/a sumffo_0/clk 0.13fF
C654 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.04fF
C655 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.04fF
C656 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.13fF
C657 ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd 0.03fF
C658 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# sumffo_0/k 0.45fF
C659 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# vdd 0.10fF
C660 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.00fF
C661 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C662 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.04fF
C663 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q 0.32fF
C664 sumffo_0/clk ffipgarr_0/y3in 0.70fF
C665 ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd 0.15fF
C666 vdd sumffo_0/ffo_0/nand_6/w_0_0# 0.10fF
C667 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C668 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 1.63fF
C669 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C670 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/x3in 0.01fF
C671 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# cla_0/g0 0.04fF
C672 vdd sumffo_0/ffo_0/d 0.04fF
C673 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C674 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.45fF
C675 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C676 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C677 ffipgarr_0/ffipg_0/ffi_1/nand_1/b vdd 0.31fF
C678 cla_1/n vdd 0.28fF
C679 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.04fF
C680 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C681 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C682 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.32fF
C683 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C684 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.31fF
C685 ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd 0.17fF
C686 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/q 0.31fF
C687 gnd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.22fF
C688 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.31fF
C689 ffipgarr_0/ffipg_2/ffi_1/qbar vdd 0.33fF
C690 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C691 cla_0/inv_0/op cla_0/nand_0/w_0_0# 0.06fF
C692 gnd sumffo_0/ffo_0/d 0.37fF
C693 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# vdd 0.10fF
C694 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# vdd 0.10fF
C695 ffipgarr_0/ffipg_2/ffi_1/inv_1/op sumffo_0/clk 0.07fF
C696 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C697 ffipgarr_0/ffipg_0/ffi_1/nand_1/b gnd 0.26fF
C698 gnd cla_1/n 0.03fF
C699 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.06fF
C700 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C701 cla_2/g0 cla_1/nor_1/w_0_0# 0.02fF
C702 ffipgarr_0/x4in ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.01fF
C703 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.06fF
C704 ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd 0.10fF
C705 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_3/b 0.33fF
C706 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# vdd 0.10fF
C707 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.04fF
C708 ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 0.13fF
C709 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C710 cla_1/g0 cla_0/inv_0/in 0.04fF
C711 ffipgarr_0/ffipg_2/ffi_1/qbar gnd 0.34fF
C712 ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd 0.34fF
C713 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C714 ffipgarr_0/ffipg_3/ffi_1/q vdd 1.35fF
C715 sumffo_0/c ffipgarr_0/ffi_0/nand_6/a 0.31fF
C716 ffipgarr_0/ffi_0/nand_6/a vdd 0.30fF
C717 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/q 0.06fF
C718 gnd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.00fF
C719 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# vdd 0.10fF
C720 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.06fF
C721 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/k3 0.46fF
C722 ffipgarr_0/ffipg_2/ffi_0/q cla_2/p0 0.03fF
C723 sumffo_0/ffo_0/inv_0/w_0_6# vdd 0.06fF
C724 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# 0.06fF
C725 ffipgarr_0/ffipg_0/ffi_0/q vdd 0.38fF
C726 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# sumffo_0/clk 0.06fF
C727 gnd cla_0/nor_1/a_13_6# 0.01fF
C728 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.33fF
C729 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.04fF
C730 ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd 0.03fF
C731 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C732 ffipgarr_0/ffipg_3/ffi_1/q gnd 0.93fF
C733 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C734 cla_2/nor_0/w_0_0# vdd 0.31fF
C735 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b 0.13fF
C736 ffipgarr_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.04fF
C737 ffipgarr_0/ffipg_3/ffi_0/q vdd 0.38fF
C738 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C739 ffipgarr_0/ffi_0/nand_6/a gnd 0.03fF
C740 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# gnd 0.00fF
C741 ffipgarr_0/ffipg_2/ffi_0/qbar vdd 0.33fF
C742 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C743 gnd ffipgarr_0/ffipg_0/ffi_0/q 2.62fF
C744 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/q 0.31fF
C745 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C746 ffipgarr_0/ffi_0/inv_1/op vdd 1.63fF
C747 sumffo_0/sbar sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C748 sumffo_0/xor_0/inv_1/op sumffo_0/k 0.06fF
C749 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C750 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/q 0.31fF
C751 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C752 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# vdd 0.10fF
C753 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# sumffo_0/clk 0.06fF
C754 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op vdd 0.15fF
C755 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C756 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C757 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.04fF
C758 ffipgarr_0/ffipg_3/ffi_0/q gnd 2.62fF
C759 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# vdd 0.10fF
C760 ffipgarr_0/ffipg_2/ffi_0/qbar gnd 0.34fF
C761 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.06fF
C762 ffipgarr_0/ffipg_3/ffi_0/nand_1/a sumffo_0/clk 0.13fF
C763 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# ffipgarr_0/x4in 0.06fF
C764 sumffo_0/c ffipgarr_0/ffi_0/nand_6/w_0_0# 0.06fF
C765 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# sumffo_0/k 0.01fF
C766 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C767 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.31fF
C768 ffipgarr_0/ffi_0/nand_6/w_0_0# vdd 0.10fF
C769 ffipgarr_0/ffi_0/inv_1/op gnd 0.22fF
C770 sumffo_0/xor_0/inv_0/op sumffo_0/c 0.20fF
C771 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C772 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# vdd 0.10fF
C773 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op vdd 0.15fF
C774 sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# 0.04fF
C775 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# gnd 0.00fF
C776 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.17fF
C777 ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd 0.34fF
C778 sumffo_0/xor_0/inv_0/op vdd 0.15fF
C779 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op vdd 0.15fF
C780 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# vdd 0.11fF
C781 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# vdd 0.11fF
C782 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C783 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C784 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C785 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C786 ffipgarr_0/k4 vdd 0.13fF
C787 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.04fF
C788 ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd 0.30fF
C789 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C790 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op gnd 0.20fF
C791 cla_0/nand_0/w_0_0# vdd 0.10fF
C792 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_1/qbar 0.06fF
C793 sumffo_0/xor_0/inv_0/op gnd 0.17fF
C794 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.17fF
C795 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# vdd 0.10fF
C796 ffipgarr_0/y2in ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.04fF
C797 ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd 0.03fF
C798 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C799 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.06fF
C800 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C801 ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 0.13fF
C802 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# sumffo_0/clk 0.06fF
C803 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.04fF
C804 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C805 ffipgarr_0/k4 gnd 0.14fF
C806 ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd 0.34fF
C807 gnd ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.14fF
C808 sumffo_0/clk ffipgarr_0/y2in 0.70fF
C809 ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd 0.30fF
C810 ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd 0.34fF
C811 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_0/q 0.73fF
C812 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C813 cla_2/p0 vdd 0.43fF
C814 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C815 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# sumffo_0/clk 0.06fF
C816 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C817 sumffo_0/c sumffo_0/xor_0/w_n3_4# 0.06fF
C818 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.06fF
C819 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C820 ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd 0.17fF
C821 cla_0/p0 cla_0/g0 0.49fF
C822 ffipgarr_0/y4in vdd 0.04fF
C823 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.04fF
C824 sumffo_0/xor_0/w_n3_4# vdd 0.12fF
C825 ffipgarr_0/x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C826 gnd ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.03fF
C827 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.04fF
C828 ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd 0.14fF
C829 gnd ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.03fF
C830 cla_2/inv_0/op vdd 0.17fF
C831 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.31fF
C832 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# vdd 0.10fF
C833 gnd cla_2/p0 0.74fF
C834 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.45fF
C835 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q 0.32fF
C836 ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd 0.34fF
C837 ffipgarr_0/ffipg_1/ffi_1/q vdd 1.35fF
C838 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# ffipgarr_0/x1in 0.06fF
C839 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q 0.32fF
C840 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.06fF
C841 ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd 0.34fF
C842 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C843 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.31fF
C844 ffipgarr_0/ffipg_1/ffi_0/q cla_1/g0 0.13fF
C845 gnd ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.10fF
C846 cla_0/nor_1/w_0_0# cla_1/g0 0.02fF
C847 ffipgarr_0/y4in gnd 0.19fF
C848 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.13fF
C849 vdd sumffo_0/ffo_0/nand_1/b 0.31fF
C850 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/w_0_0# 0.06fF
C851 cla_0/p0 vdd 0.28fF
C852 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.13fF
C853 cla_2/inv_0/op gnd 0.10fF
C854 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C855 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C856 cla_2/p1 vdd 0.31fF
C857 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q 0.32fF
C858 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# vdd 0.10fF
C859 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/q 0.31fF
C860 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# vdd 0.10fF
C861 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.31fF
C862 ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd 0.03fF
C863 ffipgarr_0/ffipg_1/ffi_1/q gnd 0.93fF
C864 ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd 0.03fF
C865 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C866 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/q 0.00fF
C867 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C868 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.13fF
C869 ffipgarr_0/x1in vdd 0.04fF
C870 ffipgarr_0/y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.04fF
C871 gnd sumffo_0/ffo_0/nand_1/b 0.26fF
C872 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# vdd 0.10fF
C873 gnd cla_0/p0 0.18fF
C874 ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 0.13fF
C875 sumffo_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C876 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.45fF
C877 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b 0.32fF
C878 ffipgarr_0/ffipg_1/ffi_1/q cla_0/p1 0.22fF
C879 gnd cla_2/p1 0.69fF
C880 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.31fF
C881 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C882 cla_1/inv_0/in cla_1/g0 0.16fF
C883 cla_0/p0 cla_0/p1 0.24fF
C884 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.13fF
C885 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.32fF
C886 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.31fF
C887 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/y4in 0.04fF
C888 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.00fF
C889 gnd ffipgarr_0/x1in 0.19fF
C890 gnd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.00fF
C891 cla_2/g0 vdd 0.47fF
C892 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# vdd 0.10fF
C893 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C894 z1o sumffo_0/ffo_0/nand_7/w_0_0# 0.04fF
C895 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C896 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# vdd 0.06fF
C897 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C898 sumffo_0/clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C899 ffipgarr_0/ffipg_2/ffi_1/q vdd 1.35fF
C900 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C901 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.06fF
C902 cla_2/g0 gnd 0.33fF
C903 ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd 0.39fF
C904 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k 0.06fF
C905 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C906 z1o sumffo_0/ffo_0/nand_6/w_0_0# 0.06fF
C907 cla_2/l vdd 0.20fF
C908 ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd 1.63fF
C909 ffipgarr_0/ffi_0/nand_5/w_0_0# vdd 0.10fF
C910 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/ffi_0/q 0.12fF
C911 cla_1/nand_0/w_0_0# vdd 0.10fF
C912 ffipgarr_0/ffipg_2/ffi_1/q gnd 0.93fF
C913 ffipgarr_0/y2in ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C914 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# vdd 0.06fF
C915 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.07fF
C916 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.32fF
C917 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C918 ffipgarr_0/ffi_0/nand_2/w_0_0# sumffo_0/clk 0.06fF
C919 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/qbar 0.31fF
C920 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_0/q 0.12fF
C921 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.06fF
C922 cla_1/l cla_1/nor_0/w_0_0# 0.05fF
C923 ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd 0.35fF
C924 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C925 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.03fF
C926 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.04fF
C927 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C928 ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd 1.63fF
C929 gnd cla_2/l 0.18fF
C930 gnd ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.22fF
C931 sumffo_0/clk sumffo_0/ffo_0/nand_0/b 0.04fF
C932 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.06fF
C933 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.33fF
C934 gnd ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# 0.01fF
C935 ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd 0.30fF
C936 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.06fF
C937 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.06fF
C938 ffipgarr_0/ffipg_3/ffi_1/qbar vdd 0.33fF
C939 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.00fF
C940 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.04fF
C941 ffipgarr_0/ffipg_0/ffi_1/qbar vdd 0.33fF
C942 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.04fF
C943 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# vdd 0.10fF
C944 ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd 0.22fF
C945 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# vdd 0.10fF
C946 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.33fF
C947 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/qbar 0.31fF
C948 sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d 0.52fF
C949 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q 0.22fF
C950 cla_2/inv_0/op cla_2/g1 0.35fF
C951 ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd 0.03fF
C952 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.31fF
C953 gnd ffipgarr_0/ffipg_3/ffi_1/qbar 0.34fF
C954 cla_1/inv_0/op vdd 0.17fF
C955 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C956 ffipgarr_0/y4in ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C957 ffipgarr_0/ffipg_0/ffi_1/qbar gnd 0.34fF
C958 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/k4 0.45fF
C959 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.03fF
C960 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C961 ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C962 ffipgarr_0/ffipg_2/ffi_1/nand_1/a sumffo_0/clk 0.13fF
C963 ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd 0.30fF
C964 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C965 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# vdd 0.11fF
C966 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_1/w_0_6# 0.03fF
C967 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# vdd 0.06fF
C968 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C969 cla_1/p0 cla_2/p0 0.24fF
C970 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# vdd 0.11fF
C971 cla_2/p1 cla_2/g1 0.00fF
C972 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.45fF
C973 gnd cla_1/inv_0/op 0.10fF
C974 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/k2 0.52fF
C975 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.04fF
C976 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.75fF
C977 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C978 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.31fF
C979 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.08fF
C980 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_0/q 0.23fF
C981 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.32fF
C982 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# sumffo_0/k 0.21fF
C983 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/k3 0.02fF
C984 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# vdd 0.11fF
C985 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# vdd 0.93fF
C986 ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd 0.14fF
C987 ffipgarr_0/cinin ffipgarr_0/ffi_0/inv_0/op 0.04fF
C988 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C989 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C990 ffipgarr_0/ffipg_1/ffi_0/nand_1/b vdd 0.31fF
C991 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b 0.13fF
C992 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/k4 0.52fF
C993 gnd cla_2/nor_1/a_13_6# 0.01fF
C994 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.04fF
C995 ffipgarr_0/ffipg_0/ffi_1/q sumffo_0/k 0.46fF
C996 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C997 cla_2/g0 cla_2/g1 0.11fF
C998 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C999 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.33fF
C1000 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.45fF
C1001 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C1002 cla_0/n vdd 0.28fF
C1003 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/k3 0.07fF
C1004 ffipgarr_0/ffipg_1/ffi_0/nand_1/b gnd 0.26fF
C1005 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b 0.13fF
C1006 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/d 0.40fF
C1007 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1008 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# cla_0/p1 0.05fF
C1009 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C1010 ffipgarr_0/cinin vdd 0.04fF
C1011 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.04fF
C1012 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# vdd 0.10fF
C1013 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C1014 cla_0/nor_0/w_0_0# vdd 0.31fF
C1015 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# cla_2/p1 0.24fF
C1016 gnd cla_0/n 0.03fF
C1017 cla_2/nor_1/w_0_0# vdd 0.31fF
C1018 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C1019 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/inv_0/op 0.06fF
C1020 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C1021 ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd 0.17fF
C1022 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# vdd 0.10fF
C1023 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.31fF
C1024 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q 0.22fF
C1025 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.31fF
C1026 ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd 0.30fF
C1027 ffipgarr_0/cinin gnd 0.19fF
C1028 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.06fF
C1029 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q 0.27fF
C1030 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.04fF
C1031 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.04fF
C1032 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C1033 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1034 ffipgarr_0/k2 ffipgarr_0/ffipg_1/ffi_1/q 0.46fF
C1035 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1036 cla_2/nor_1/w_0_0# gnd 0.01fF
C1037 ffipgarr_0/ffi_0/inv_1/w_0_6# sumffo_0/clk 0.06fF
C1038 vdd sumffo_0/ffo_0/inv_0/op 0.17fF
C1039 sumffo_0/clk ffipgarr_0/x2in 0.70fF
C1040 ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd 0.39fF
C1041 gnd ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.10fF
C1042 ffipgarr_0/k2 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C1043 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C1044 ffipgarr_0/x4in vdd 0.04fF
C1045 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.31fF
C1046 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.00fF
C1047 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C1048 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.04fF
C1049 cla_0/p1 cla_0/nor_0/w_0_0# 0.06fF
C1050 ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd 0.03fF
C1051 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C1052 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# vdd 0.10fF
C1053 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# vdd 0.10fF
C1054 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# vdd 0.11fF
C1055 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.03fF
C1056 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/q 0.31fF
C1057 gnd sumffo_0/ffo_0/inv_0/op 0.10fF
C1058 ffipgarr_0/x3in sumffo_0/clk 0.70fF
C1059 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.13fF
C1060 ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd 0.35fF
C1061 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C1062 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C1063 ffipgarr_0/x4in gnd 0.19fF
C1064 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# vdd 0.06fF
C1065 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/k3 0.45fF
C1066 cla_1/nor_1/w_0_0# vdd 0.31fF
C1067 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# vdd 0.06fF
C1068 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.32fF
C1069 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.32fF
C1070 ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd 0.39fF
C1071 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.04fF
C1072 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C1073 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# vdd 0.10fF
C1074 ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd 0.30fF
C1075 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/cinbar 0.31fF
C1076 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.04fF
C1077 sumffo_0/ffo_0/nand_1/a vdd 0.30fF
C1078 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.04fF
C1079 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C1080 vdd sumffo_0/ffo_0/nand_3/w_0_0# 0.11fF
C1081 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op vdd 0.15fF
C1082 gnd cla_1/nor_1/w_0_0# 0.01fF
C1083 ffipgarr_0/k3 vdd 0.13fF
C1084 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1085 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_0/q 0.73fF
C1086 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C1087 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C1088 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# vdd 0.10fF
C1089 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/w_n3_4# 0.06fF
C1090 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/qbar 0.00fF
C1091 ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd 1.63fF
C1092 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.03fF
C1093 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.35fF
C1094 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1095 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# vdd 0.10fF
C1096 gnd ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.03fF
C1097 cla_1/inv_0/in cla_2/p0 0.02fF
C1098 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.04fF
C1099 sumffo_0/ffo_0/nand_1/a gnd 0.03fF
C1100 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# sumffo_0/clk 0.06fF
C1101 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a 0.00fF
C1102 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C1103 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C1104 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# cla_2/p0 0.24fF
C1105 ffipgarr_0/k3 gnd 0.14fF
C1106 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/w_0_0# 0.06fF
C1107 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# vdd 0.11fF
C1108 ffipgarr_0/ffipg_0/ffi_0/q sumffo_0/k 0.07fF
C1109 ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd 0.22fF
C1110 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.32fF
C1111 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.04fF
C1112 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C1113 ffipgarr_0/ffipg_1/ffi_1/nand_1/b vdd 0.31fF
C1114 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.33fF
C1115 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.04fF
C1116 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/k4 0.21fF
C1117 ffipgarr_0/ffi_0/inv_0/w_0_6# ffipgarr_0/cinin 0.06fF
C1118 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.31fF
C1119 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C1120 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C1121 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# 0.04fF
C1122 sumffo_0/clk sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1123 sumffo_0/clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.13fF
C1124 ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd 0.30fF
C1125 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C1126 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_1/b 0.45fF
C1127 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.13fF
C1128 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# vdd 0.06fF
C1129 ffipgarr_0/x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.04fF
C1130 ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd 1.63fF
C1131 ffipgarr_0/x4in ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.04fF
C1132 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C1133 ffipgarr_0/ffi_0/nand_4/w_0_0# vdd 0.10fF
C1134 ffipgarr_0/ffipg_1/ffi_1/nand_1/b gnd 0.26fF
C1135 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/q 0.31fF
C1136 sumffo_0/clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.13fF
C1137 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# vdd 0.10fF
C1138 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.04fF
C1139 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.32fF
C1140 cla_2/nor_1/w_0_0# cla_2/g1 0.02fF
C1141 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C1142 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.03fF
C1143 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_0/q 0.12fF
C1144 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.04fF
C1145 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/q 0.20fF
C1146 cla_0/inv_0/op vdd 0.17fF
C1147 ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd 0.22fF
C1148 vdd sumffo_0/ffo_0/nand_2/w_0_0# 0.10fF
C1149 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# vdd 0.10fF
C1150 sumffo_0/xor_0/inv_0/op sumffo_0/k 0.27fF
C1151 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C1152 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C1153 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.04fF
C1154 sumffo_0/clk ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.07fF
C1155 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.04fF
C1156 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C1157 sumffo_0/c sumffo_0/xor_0/a_10_10# 0.12fF
C1158 sumffo_0/clk sumffo_0/ffo_0/d 0.04fF
C1159 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.04fF
C1160 ffipgarr_0/ffipg_2/ffi_0/q vdd 0.38fF
C1161 gnd cla_0/inv_0/op 0.10fF
C1162 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.06fF
C1163 cla_2/g0 cla_1/inv_0/in 0.04fF
C1164 vdd sumffo_0/xor_0/a_10_10# 0.93fF
C1165 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.06fF
C1166 sumffo_0/ffo_0/nand_5/w_0_0# vdd 0.10fF
C1167 ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd 0.30fF
C1168 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.04fF
C1169 ffipgarr_0/cinbar ffipgarr_0/ffi_0/nand_6/a 0.00fF
C1170 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C1171 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# cla_2/g0 0.04fF
C1172 sumffo_0/clk ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.32fF
C1173 cla_1/l cla_2/p0 0.02fF
C1174 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1175 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1176 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1177 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1178 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1179 sumffo_0/k Gnd 3.91fF
C1180 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1181 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1182 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1183 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1184 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1185 sumffo_0/sbar Gnd 0.43fF
C1186 vdd Gnd 19.28fF
C1187 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1188 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1189 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1190 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1191 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1192 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1193 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1194 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1195 sumffo_0/ffo_0/d Gnd 0.64fF
C1196 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1197 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1198 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1199 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1200 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1201 cla_2/p1 Gnd 1.09fF
C1202 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1203 cla_2/l Gnd 0.06fF
C1204 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1205 cla_2/inv_0/in Gnd 0.27fF
C1206 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1207 gnd Gnd 32.63fF
C1208 cla_2/n Gnd 0.09fF
C1209 cla_2/g1 Gnd 0.60fF
C1210 cla_2/inv_0/op Gnd 0.26fF
C1211 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1212 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1213 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1214 ffipgarr_0/ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1215 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1216 ffipgarr_0/ffipg_3/ffi_1/qbar Gnd 0.42fF
C1217 ffipgarr_0/ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1218 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1219 ffipgarr_0/ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1220 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1221 ffipgarr_0/ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1222 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1223 ffipgarr_0/ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1224 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1225 ffipgarr_0/x4in Gnd 0.51fF
C1226 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1227 ffipgarr_0/ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1228 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1229 ffipgarr_0/ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1230 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1231 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1232 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1233 ffipgarr_0/ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1234 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1235 ffipgarr_0/ffipg_3/ffi_0/qbar Gnd 0.42fF
C1236 ffipgarr_0/ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1237 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1238 ffipgarr_0/ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1239 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1240 ffipgarr_0/ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1241 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1242 ffipgarr_0/ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1243 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1244 ffipgarr_0/y4in Gnd 0.51fF
C1245 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1246 ffipgarr_0/ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1247 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1248 ffipgarr_0/ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C1249 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1250 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1251 ffipgarr_0/k4 Gnd 1.10fF
C1252 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1253 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1254 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1255 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1256 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1257 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1258 ffipgarr_0/ffipg_3/ffi_0/q Gnd 2.68fF
C1259 ffipgarr_0/ffipg_3/ffi_1/q Gnd 2.93fF
C1260 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1261 ffipgarr_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1262 ffipgarr_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1263 sumffo_0/c Gnd 1.70fF
C1264 ffipgarr_0/ffi_0/nand_7/a Gnd 0.30fF
C1265 ffipgarr_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1266 ffipgarr_0/cinbar Gnd 0.44fF
C1267 ffipgarr_0/ffi_0/nand_6/a Gnd 0.30fF
C1268 ffipgarr_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1269 ffipgarr_0/ffi_0/inv_1/op Gnd 0.89fF
C1270 ffipgarr_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1271 ffipgarr_0/ffi_0/nand_3/b Gnd 0.43fF
C1272 ffipgarr_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1273 ffipgarr_0/ffi_0/nand_3/a Gnd 0.30fF
C1274 ffipgarr_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1275 sumffo_0/clk Gnd 13.01fF
C1276 ffipgarr_0/cinin Gnd 0.50fF
C1277 ffipgarr_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1278 ffipgarr_0/ffi_0/inv_0/op Gnd 0.26fF
C1279 ffipgarr_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1280 ffipgarr_0/ffi_0/nand_1/a Gnd 0.30fF
C1281 ffipgarr_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1282 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1283 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1284 ffipgarr_0/ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C1285 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1286 ffipgarr_0/ffipg_2/ffi_1/qbar Gnd 0.42fF
C1287 ffipgarr_0/ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C1288 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1289 ffipgarr_0/ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C1290 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1291 ffipgarr_0/ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C1292 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1293 ffipgarr_0/ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C1294 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1295 ffipgarr_0/x3in Gnd 0.51fF
C1296 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1297 ffipgarr_0/ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C1298 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1299 ffipgarr_0/ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C1300 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1301 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1302 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1303 ffipgarr_0/ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C1304 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1305 ffipgarr_0/ffipg_2/ffi_0/qbar Gnd 0.42fF
C1306 ffipgarr_0/ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C1307 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1308 ffipgarr_0/ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C1309 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1310 ffipgarr_0/ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C1311 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1312 ffipgarr_0/ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C1313 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1314 ffipgarr_0/y3in Gnd 0.51fF
C1315 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1316 ffipgarr_0/ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C1317 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1318 ffipgarr_0/ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C1319 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1320 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1321 ffipgarr_0/k3 Gnd 1.10fF
C1322 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1323 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1324 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1325 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1326 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1327 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1328 ffipgarr_0/ffipg_2/ffi_0/q Gnd 2.68fF
C1329 ffipgarr_0/ffipg_2/ffi_1/q Gnd 2.93fF
C1330 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1331 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1332 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1333 ffipgarr_0/ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C1334 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1335 ffipgarr_0/ffipg_1/ffi_1/qbar Gnd 0.42fF
C1336 ffipgarr_0/ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C1337 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1338 ffipgarr_0/ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C1339 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1340 ffipgarr_0/ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C1341 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1342 ffipgarr_0/ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C1343 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1344 ffipgarr_0/x2in Gnd 0.51fF
C1345 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1346 ffipgarr_0/ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C1347 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1348 ffipgarr_0/ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C1349 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1350 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1351 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1352 ffipgarr_0/ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C1353 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1354 ffipgarr_0/ffipg_1/ffi_0/qbar Gnd 0.42fF
C1355 ffipgarr_0/ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C1356 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1357 ffipgarr_0/ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C1358 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1359 ffipgarr_0/ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C1360 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1361 ffipgarr_0/ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C1362 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1363 ffipgarr_0/y2in Gnd 0.51fF
C1364 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1365 ffipgarr_0/ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C1366 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1367 ffipgarr_0/ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C1368 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1369 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1370 ffipgarr_0/k2 Gnd 1.10fF
C1371 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1372 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1373 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1374 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1375 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1376 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1377 ffipgarr_0/ffipg_1/ffi_0/q Gnd 2.68fF
C1378 ffipgarr_0/ffipg_1/ffi_1/q Gnd 2.93fF
C1379 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1380 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1381 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1382 ffipgarr_0/ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C1383 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1384 ffipgarr_0/ffipg_0/ffi_1/qbar Gnd 0.42fF
C1385 ffipgarr_0/ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C1386 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1387 ffipgarr_0/ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C1388 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1389 ffipgarr_0/ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C1390 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1391 ffipgarr_0/ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C1392 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1393 ffipgarr_0/x1in Gnd 0.51fF
C1394 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1395 ffipgarr_0/ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C1396 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1397 ffipgarr_0/ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C1398 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1399 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1400 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1401 ffipgarr_0/ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C1402 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1403 ffipgarr_0/ffipg_0/ffi_0/qbar Gnd 0.42fF
C1404 ffipgarr_0/ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C1405 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1406 ffipgarr_0/ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C1407 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1408 ffipgarr_0/ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C1409 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1410 ffipgarr_0/ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C1411 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1412 ffipgarr_0/y1in Gnd 0.51fF
C1413 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1414 ffipgarr_0/ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C1415 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1416 ffipgarr_0/ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C1417 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1418 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1419 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1420 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1421 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1422 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1423 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1424 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1425 cla_0/g0 Gnd 1.41fF
C1426 ffipgarr_0/ffipg_0/ffi_0/q Gnd 2.68fF
C1427 ffipgarr_0/ffipg_0/ffi_1/q Gnd 2.93fF
C1428 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1429 cla_2/p0 Gnd 1.75fF
C1430 cla_1/nor_1/w_0_0# Gnd 1.23fF
C1431 cla_1/l Gnd 0.06fF
C1432 cla_1/p0 Gnd 0.20fF
C1433 cla_1/nor_0/w_0_0# Gnd 1.23fF
C1434 cla_1/inv_0/in Gnd 0.27fF
C1435 cla_1/inv_0/w_0_6# Gnd 0.58fF
C1436 cla_1/n Gnd 0.09fF
C1437 cla_1/inv_0/op Gnd 0.26fF
C1438 cla_1/nand_0/w_0_0# Gnd 0.82fF
C1439 cla_0/p1 Gnd 1.59fF
C1440 cla_0/nor_1/w_0_0# Gnd 1.23fF
C1441 cla_0/l Gnd 0.06fF
C1442 cla_0/nor_0/w_0_0# Gnd 1.23fF
C1443 cla_0/inv_0/in Gnd 0.27fF
C1444 cla_0/inv_0/w_0_6# Gnd 0.58fF
C1445 cla_0/n Gnd 0.09fF
C1446 cla_1/g0 Gnd 0.85fF
C1447 cla_0/inv_0/op Gnd 0.26fF
C1448 cla_0/nand_0/w_0_0# Gnd 0.82fF
