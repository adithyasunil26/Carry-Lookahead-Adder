magic
tech scmos
timestamp 1618536408
<< nwell >>
rect 0 6 24 30
<< polysilicon >>
rect 11 24 13 27
rect 11 -2 13 12
rect 11 -11 13 -8
<< ndiffusion >>
rect 6 -4 11 -2
rect 10 -8 11 -4
rect 13 -6 14 -2
rect 13 -8 18 -6
<< pdiffusion >>
rect 10 20 11 24
rect 6 12 11 20
rect 13 16 18 24
rect 13 12 14 16
<< metal1 >>
rect 0 30 24 33
rect 6 24 9 30
rect 15 5 18 12
rect 0 2 7 5
rect 15 2 24 5
rect 15 -2 18 2
rect 6 -12 9 -8
rect 0 -15 24 -12
<< ntransistor >>
rect 11 -8 13 -2
<< ptransistor >>
rect 11 12 13 24
<< polycontact >>
rect 7 1 11 5
<< ndcontact >>
rect 6 -8 10 -4
rect 14 -6 18 -2
<< pdcontact >>
rect 6 20 10 24
rect 14 12 18 16
<< labels >>
rlabel metal1 14 31 14 31 5 vdd!
rlabel metal1 24 2 24 5 7 op
rlabel metal1 0 2 0 5 3 in
rlabel metal1 20 -14 20 -14 1 gnd!
<< end >>
