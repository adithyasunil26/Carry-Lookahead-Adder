* SPICE3 file created from ckt.ext - technology: scmos

.option scale=0.09u

M1000 ffipg_6/pggen_0/nand_0/a_13_n26# ffipg_6/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=17130 ps=10312
M1001 gnd ffipg_6/ffi_0/q ffipg_6/g ffipg_6/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=34260 pd=18984 as=96 ps=40
M1002 ffipg_6/g ffipg_6/ffi_1/q gnd ffipg_6/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 ffipg_6/g ffipg_6/ffi_0/q ffipg_6/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1005 ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/ffi_1/q gnd ffipg_6/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1006 ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1007 ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/ffi_0/q gnd ffipg_6/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 gnd ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/a_10_10# ffipg_6/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1009 ffipg_6/k ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1010 gnd ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1011 ffipg_6/pggen_0/xor_0/a_10_10# ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/k ffipg_6/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1012 ffipg_6/pggen_0/xor_0/a_10_n43# ffipg_6/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 ffipg_6/pggen_0/xor_0/a_38_n43# ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 ffipg_6/pggen_0/xor_0/a_10_10# ffipg_6/ffi_1/q gnd ffipg_6/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 ffipg_6/k ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/pggen_0/xor_0/a_10_10# ffipg_6/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 ffipg_6/p ffipg_6/ffi_1/q ffipg_6/pggen_0/nor_0/a_13_6# ffipg_6/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1017 ffipg_6/pggen_0/nor_0/a_13_6# ffipg_6/ffi_0/q gnd ffipg_6/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 gnd ffipg_6/ffi_1/q ffipg_6/p Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1019 ffipg_6/p ffipg_6/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 ffipg_6/ffi_0/nand_1/a_13_n26# ffipg_6/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_1/a gnd ffipg_6/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 ffipg_6/ffi_0/nand_0/a_13_n26# ffipg_6/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1025 gnd clk ffipg_6/ffi_0/nand_1/a ffipg_6/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1026 ffipg_6/ffi_0/nand_1/a ffipg_6/ffi_0/inv_0/op gnd ffipg_6/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 ffipg_6/ffi_0/nand_1/a clk ffipg_6/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1028 ffipg_6/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1029 gnd clk ffipg_6/ffi_0/nand_3/a ffipg_6/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1030 ffipg_6/ffi_0/nand_3/a y3in gnd ffipg_6/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 ffipg_6/ffi_0/nand_3/a clk ffipg_6/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1032 ffipg_6/ffi_0/nand_3/a_13_n26# ffipg_6/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1033 gnd ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1034 ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_3/a gnd ffipg_6/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1036 ffipg_6/ffi_0/nand_4/a_13_n26# ffipg_6/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1037 gnd ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_0/nand_6/a ffipg_6/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1038 ffipg_6/ffi_0/nand_6/a ffipg_6/ffi_0/nand_3/b gnd ffipg_6/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 ffipg_6/ffi_0/nand_6/a ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1040 ffipg_6/ffi_0/nand_5/a_13_n26# ffipg_6/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1041 gnd ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_7/a ffipg_6/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1042 ffipg_6/ffi_0/nand_7/a ffipg_6/ffi_0/inv_1/op gnd ffipg_6/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 ffipg_6/ffi_0/nand_7/a ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 ffipg_6/ffi_0/nand_6/a_13_n26# ffipg_6/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1045 gnd ffipg_6/ffi_0/q ffipg_6/ffi_0/qbar ffipg_6/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1046 ffipg_6/ffi_0/qbar ffipg_6/ffi_0/nand_6/a gnd ffipg_6/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 ffipg_6/ffi_0/qbar ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1048 ffipg_6/ffi_0/nand_7/a_13_n26# ffipg_6/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1049 gnd ffipg_6/ffi_0/qbar ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1050 ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_7/a gnd ffipg_6/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 ffipg_6/ffi_0/q ffipg_6/ffi_0/qbar ffipg_6/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1052 ffipg_6/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1053 ffipg_6/ffi_0/inv_0/op y3in gnd ffipg_6/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1054 ffipg_6/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1055 ffipg_6/ffi_0/inv_1/op clk gnd ffipg_6/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 ffipg_6/ffi_1/nand_1/a_13_n26# ffipg_6/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1057 gnd ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/b ffipg_6/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1058 ffipg_6/ffi_1/nand_3/b ffipg_6/ffi_1/nand_1/a gnd ffipg_6/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 ffipg_6/ffi_1/nand_3/b ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1060 ffipg_6/ffi_1/nand_0/a_13_n26# ffipg_6/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1061 gnd clk ffipg_6/ffi_1/nand_1/a ffipg_6/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1062 ffipg_6/ffi_1/nand_1/a ffipg_6/ffi_1/inv_0/op gnd ffipg_6/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 ffipg_6/ffi_1/nand_1/a clk ffipg_6/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1064 ffipg_6/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1065 gnd clk ffipg_6/ffi_1/nand_3/a ffipg_6/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1066 ffipg_6/ffi_1/nand_3/a x3in gnd ffipg_6/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 ffipg_6/ffi_1/nand_3/a clk ffipg_6/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 ffipg_6/ffi_1/nand_3/a_13_n26# ffipg_6/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1069 gnd ffipg_6/ffi_1/nand_3/b ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1070 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/a gnd ffipg_6/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/b ffipg_6/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1072 ffipg_6/ffi_1/nand_4/a_13_n26# ffipg_6/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1073 gnd ffipg_6/ffi_1/inv_1/op ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1074 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/nand_3/b gnd ffipg_6/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/inv_1/op ffipg_6/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1076 ffipg_6/ffi_1/nand_5/a_13_n26# ffipg_6/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1077 gnd ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_7/a ffipg_6/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1078 ffipg_6/ffi_1/nand_7/a ffipg_6/ffi_1/inv_1/op gnd ffipg_6/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 ffipg_6/ffi_1/nand_7/a ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 ffipg_6/ffi_1/nand_6/a_13_n26# ffipg_6/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1081 gnd ffipg_6/ffi_1/q ffipg_6/ffi_1/qbar ffipg_6/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1082 ffipg_6/ffi_1/qbar ffipg_6/ffi_1/nand_6/a gnd ffipg_6/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 ffipg_6/ffi_1/qbar ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1084 ffipg_6/ffi_1/nand_7/a_13_n26# ffipg_6/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 gnd ffipg_6/ffi_1/qbar ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1086 ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_7/a gnd ffipg_6/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 ffipg_6/ffi_1/q ffipg_6/ffi_1/qbar ffipg_6/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1088 ffipg_6/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1089 ffipg_6/ffi_1/inv_0/op x3in gnd ffipg_6/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1090 ffipg_6/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 ffipg_6/ffi_1/inv_1/op clk gnd ffipg_6/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 ffipg_7/pggen_0/nand_0/a_13_n26# ffipg_7/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 gnd ffipg_7/ffi_0/q ffipg_7/g ffipg_7/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1094 ffipg_7/g ffipg_7/ffi_1/q gnd ffipg_7/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 ffipg_7/g ffipg_7/ffi_0/q ffipg_7/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1096 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1097 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/ffi_1/q gnd ffipg_7/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1098 ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1099 ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/ffi_0/q gnd ffipg_7/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 gnd ffipg_7/ffi_0/q ffipg_7/pggen_0/xor_0/a_10_10# ffipg_7/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1101 ffipg_7/k ffipg_7/ffi_0/q ffipg_7/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1102 gnd ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1103 ffipg_7/pggen_0/xor_0/a_10_10# ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/k ffipg_7/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1104 ffipg_7/pggen_0/xor_0/a_10_n43# ffipg_7/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 ffipg_7/pggen_0/xor_0/a_38_n43# ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 ffipg_7/pggen_0/xor_0/a_10_10# ffipg_7/ffi_1/q gnd ffipg_7/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 ffipg_7/k ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/pggen_0/xor_0/a_10_10# ffipg_7/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 ffipg_7/p ffipg_7/ffi_1/q ffipg_7/pggen_0/nor_0/a_13_6# ffipg_7/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1109 ffipg_7/pggen_0/nor_0/a_13_6# ffipg_7/ffi_0/q gnd ffipg_7/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 gnd ffipg_7/ffi_1/q ffipg_7/p Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1111 ffipg_7/p ffipg_7/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 ffipg_7/ffi_0/nand_1/a_13_n26# ffipg_7/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1113 gnd ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1114 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/a gnd ffipg_7/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 ffipg_7/ffi_0/nand_0/a_13_n26# ffipg_7/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1117 gnd clk ffipg_7/ffi_0/nand_1/a ffipg_7/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1118 ffipg_7/ffi_0/nand_1/a ffipg_7/ffi_0/inv_0/op gnd ffipg_7/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 ffipg_7/ffi_0/nand_1/a clk ffipg_7/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 ffipg_7/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 gnd clk ffipg_7/ffi_0/nand_3/a ffipg_7/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1122 ffipg_7/ffi_0/nand_3/a y4in gnd ffipg_7/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 ffipg_7/ffi_0/nand_3/a clk ffipg_7/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1124 ffipg_7/ffi_0/nand_3/a_13_n26# ffipg_7/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1125 gnd ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1126 ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_3/a gnd ffipg_7/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1128 ffipg_7/ffi_0/nand_4/a_13_n26# ffipg_7/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1129 gnd ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_0/nand_6/a ffipg_7/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1130 ffipg_7/ffi_0/nand_6/a ffipg_7/ffi_0/nand_3/b gnd ffipg_7/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 ffipg_7/ffi_0/nand_6/a ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 ffipg_7/ffi_0/nand_5/a_13_n26# ffipg_7/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1133 gnd ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_7/a ffipg_7/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1134 ffipg_7/ffi_0/nand_7/a ffipg_7/ffi_0/inv_1/op gnd ffipg_7/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ffipg_7/ffi_0/nand_7/a ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1136 ffipg_7/ffi_0/nand_6/a_13_n26# ffipg_7/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1137 gnd ffipg_7/ffi_0/q ffipg_7/ffi_0/qbar ffipg_7/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1138 ffipg_7/ffi_0/qbar ffipg_7/ffi_0/nand_6/a gnd ffipg_7/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 ffipg_7/ffi_0/qbar ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1140 ffipg_7/ffi_0/nand_7/a_13_n26# ffipg_7/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1141 gnd ffipg_7/ffi_0/qbar ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1142 ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_7/a gnd ffipg_7/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 ffipg_7/ffi_0/q ffipg_7/ffi_0/qbar ffipg_7/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 ffipg_7/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1145 ffipg_7/ffi_0/inv_0/op y4in gnd ffipg_7/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1146 ffipg_7/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1147 ffipg_7/ffi_0/inv_1/op clk gnd ffipg_7/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 ffipg_7/ffi_1/nand_1/a_13_n26# ffipg_7/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1149 gnd ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1150 ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_1/a gnd ffipg_7/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_7/ffi_1/nand_0/a_13_n26# ffipg_7/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 gnd clk ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/inv_0/op gnd ffipg_7/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 ffipg_7/ffi_1/nand_1/a clk ffipg_7/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_7/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1157 gnd clk ffipg_7/ffi_1/nand_3/a ffipg_7/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1158 ffipg_7/ffi_1/nand_3/a x4in gnd ffipg_7/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 ffipg_7/ffi_1/nand_3/a clk ffipg_7/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 ffipg_7/ffi_1/nand_3/a_13_n26# ffipg_7/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1161 gnd ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1162 ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_3/a gnd ffipg_7/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1163 ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1164 ffipg_7/ffi_1/nand_4/a_13_n26# ffipg_7/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1165 gnd ffipg_7/ffi_1/inv_1/op ffipg_7/ffi_1/nand_6/a ffipg_7/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1166 ffipg_7/ffi_1/nand_6/a ffipg_7/ffi_1/nand_3/b gnd ffipg_7/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_7/ffi_1/nand_6/a ffipg_7/ffi_1/inv_1/op ffipg_7/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1168 ffipg_7/ffi_1/nand_5/a_13_n26# ffipg_7/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1169 gnd ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_7/a ffipg_7/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1170 ffipg_7/ffi_1/nand_7/a ffipg_7/ffi_1/inv_1/op gnd ffipg_7/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ffipg_7/ffi_1/nand_7/a ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1172 ffipg_7/ffi_1/nand_6/a_13_n26# ffipg_7/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1173 gnd ffipg_7/ffi_1/q ffipg_7/ffi_1/qbar ffipg_7/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1174 ffipg_7/ffi_1/qbar ffipg_7/ffi_1/nand_6/a gnd ffipg_7/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 ffipg_7/ffi_1/qbar ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1176 ffipg_7/ffi_1/nand_7/a_13_n26# ffipg_7/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1177 gnd ffipg_7/ffi_1/qbar ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1178 ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_7/a gnd ffipg_7/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 ffipg_7/ffi_1/q ffipg_7/ffi_1/qbar ffipg_7/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_7/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_7/ffi_1/inv_0/op x4in gnd ffipg_7/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 ffipg_7/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1183 ffipg_7/ffi_1/inv_1/op clk gnd ffipg_7/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1184 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1185 gnd ffi_0/q inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1186 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 inv_2/in ffi_0/q nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1188 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1189 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1190 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1192 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1193 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1194 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1197 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1198 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1201 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1202 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1204 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1205 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1206 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1208 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1209 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1210 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1211 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1213 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1215 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1217 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1219 gnd ffi_0/q inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1220 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 inv_8/in ffi_0/q nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1223 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1224 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1226 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1227 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1228 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1229 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1231 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1233 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1235 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1237 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1238 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1240 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1241 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1243 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1245 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1247 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1249 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1251 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1252 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a gnd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1253 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1254 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1255 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1256 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op gnd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1258 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1259 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1260 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1262 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1263 gnd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1264 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a gnd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1266 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1267 gnd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1268 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b gnd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1270 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1271 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1272 sumffo_0/ffo_0/nand_7/a clk gnd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1274 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1275 gnd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1276 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a gnd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1278 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1279 gnd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1280 z1o sumffo_0/ffo_0/nand_7/a gnd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1282 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1283 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1284 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1285 sumffo_0/ffo_0/nand_0/b clk gnd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1286 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1287 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1288 sumffo_0/xor_0/inv_1/op ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1289 sumffo_0/xor_0/inv_1/op ffi_0/q gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 gnd ffi_0/q sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1291 sumffo_0/ffo_0/d ffi_0/q sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1292 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1293 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1294 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1296 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1299 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1300 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a gnd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1302 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1303 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1304 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op gnd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1305 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1306 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1307 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1308 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1309 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1310 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1311 gnd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1312 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a gnd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1313 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1314 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1315 gnd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1316 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b gnd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1317 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1318 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1319 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1320 sumffo_2/ffo_0/nand_7/a clk gnd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1321 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1322 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1323 gnd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1324 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a gnd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1325 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1326 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1327 gnd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1328 z3o sumffo_2/ffo_0/nand_7/a gnd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1330 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1331 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1333 sumffo_2/ffo_0/nand_0/b clk gnd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1334 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1335 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1337 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1338 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1339 sumffo_2/ffo_0/d ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1340 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1341 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1342 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1347 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1348 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a gnd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1350 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1351 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1352 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op gnd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1353 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1354 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1355 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1356 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1358 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1359 gnd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1360 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a gnd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1361 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1362 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1363 gnd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1364 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b gnd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1366 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1367 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1368 sumffo_1/ffo_0/nand_7/a clk gnd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1370 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1371 gnd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1372 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a gnd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1373 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1374 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1375 gnd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1376 z2o sumffo_1/ffo_0/nand_7/a gnd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1378 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1379 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1380 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1381 sumffo_1/ffo_0/nand_0/b clk gnd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1382 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1383 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1384 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1385 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1386 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1387 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1388 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1389 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1390 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1393 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1395 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1396 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a gnd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1397 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1398 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1399 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1400 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op gnd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1401 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1402 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1403 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1404 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1406 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1407 gnd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1408 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a gnd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1410 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1411 gnd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1412 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b gnd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1413 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1414 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1415 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1416 sumffo_3/ffo_0/nand_7/a clk gnd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1418 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1419 gnd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1420 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a gnd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1421 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1422 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1423 gnd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1424 z4o sumffo_3/ffo_0/nand_7/a gnd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1425 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1426 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1427 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1428 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1429 sumffo_3/ffo_0/nand_0/b clk gnd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1430 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1431 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1433 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1434 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1435 sumffo_3/ffo_0/d ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1436 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1437 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1438 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1443 gnd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1444 ffo_0/nand_3/b ffo_0/nand_1/a gnd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1445 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1446 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1447 gnd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1448 ffo_0/nand_1/a ffo_0/inv_0/op gnd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1450 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1451 gnd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1452 ffo_0/nand_3/a ffo_0/d gnd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1455 gnd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1456 ffo_0/nand_1/b ffo_0/nand_3/a gnd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1458 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1459 gnd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1460 ffo_0/nand_6/a ffo_0/nand_3/b gnd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1463 gnd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1464 ffo_0/nand_7/a clk gnd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1466 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1467 gnd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1468 ffo_0/qbar ffo_0/nand_6/a gnd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1470 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 gnd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 couto ffo_0/nand_7/a gnd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1475 ffo_0/inv_0/op ffo_0/d gnd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1476 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1477 ffo_0/nand_0/b clk gnd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1480 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1481 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1483 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1484 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1485 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1486 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1487 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1489 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1491 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1493 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1495 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1496 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1497 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1499 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1500 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1501 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1503 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1504 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1505 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1507 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1508 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1509 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1511 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1512 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1513 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1514 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1515 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1516 ffipg_0/pggen_0/nand_0/a_13_n26# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1517 gnd ffipg_0/ffi_0/q cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1518 cla_0/g0 ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1519 cla_0/g0 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1520 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1521 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1522 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1523 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1524 gnd ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1525 ffipg_0/k ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1526 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1527 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1528 ffipg_0/pggen_0/xor_0/a_10_n43# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1529 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 nor_0/a ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1533 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1534 gnd ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1535 nor_0/a ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 ffipg_0/ffi_0/nand_1/a_13_n26# ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1537 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1538 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/a gnd ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1539 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1540 ffipg_0/ffi_0/nand_0/a_13_n26# ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1541 gnd clk ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1542 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/inv_0/op gnd ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1543 ffipg_0/ffi_0/nand_1/a clk ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1544 ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1545 gnd clk ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1546 ffipg_0/ffi_0/nand_3/a y1in gnd ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1547 ffipg_0/ffi_0/nand_3/a clk ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1548 ffipg_0/ffi_0/nand_3/a_13_n26# ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1549 gnd ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1550 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/a gnd ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1551 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1552 ffipg_0/ffi_0/nand_4/a_13_n26# ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1553 gnd ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1554 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_3/b gnd ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1555 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1556 ffipg_0/ffi_0/nand_5/a_13_n26# ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1557 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1558 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/inv_1/op gnd ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1560 ffipg_0/ffi_0/nand_6/a_13_n26# ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1561 gnd ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1562 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/a gnd ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1564 ffipg_0/ffi_0/nand_7/a_13_n26# ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1565 gnd ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1566 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a gnd ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1567 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1568 ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1569 ffipg_0/ffi_0/inv_0/op y1in gnd ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1571 ffipg_0/ffi_0/inv_1/op clk gnd ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1572 ffipg_0/ffi_1/nand_1/a_13_n26# ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1573 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1574 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a gnd ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1575 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1576 ffipg_0/ffi_1/nand_0/a_13_n26# ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1577 gnd clk ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1578 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/inv_0/op gnd ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1579 ffipg_0/ffi_1/nand_1/a clk ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1580 ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1581 gnd clk ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1582 ffipg_0/ffi_1/nand_3/a x1in gnd ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1583 ffipg_0/ffi_1/nand_3/a clk ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1584 ffipg_0/ffi_1/nand_3/a_13_n26# ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1585 gnd ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1586 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/a gnd ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1587 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1588 ffipg_0/ffi_1/nand_4/a_13_n26# ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1589 gnd ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1590 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_3/b gnd ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1592 ffipg_0/ffi_1/nand_5/a_13_n26# ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1593 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1594 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/inv_1/op gnd ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1595 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1596 ffipg_0/ffi_1/nand_6/a_13_n26# ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1597 gnd ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1598 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/a gnd ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1599 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1600 ffipg_0/ffi_1/nand_7/a_13_n26# ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1601 gnd ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1602 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a gnd ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1603 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1604 ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1605 ffipg_0/ffi_1/inv_0/op x1in gnd ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1607 ffipg_0/ffi_1/inv_1/op clk gnd ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1608 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1609 ffo_0/d inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1610 ffipg_1/pggen_0/nand_0/a_13_n26# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1611 gnd ffipg_1/ffi_0/q cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 cla_0/l ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 cla_0/l ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1614 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1615 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1616 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1617 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 gnd ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1619 ffipg_1/k ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1620 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1621 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1622 ffipg_1/pggen_0/xor_0/a_10_n43# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1623 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1626 cla_1/p0 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1627 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1628 gnd ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1629 cla_1/p0 ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1630 ffipg_1/ffi_0/nand_1/a_13_n26# ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a gnd ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 ffipg_1/ffi_0/nand_0/a_13_n26# ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 gnd clk ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/inv_0/op gnd ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 ffipg_1/ffi_0/nand_1/a clk ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 gnd clk ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 ffipg_1/ffi_0/nand_3/a y2in gnd ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 ffipg_1/ffi_0/nand_3/a clk ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 ffipg_1/ffi_0/nand_3/a_13_n26# ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1643 gnd ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1644 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/a gnd ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1645 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 ffipg_1/ffi_0/nand_4/a_13_n26# ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1647 gnd ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1648 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_3/b gnd ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1649 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 ffipg_1/ffi_0/nand_5/a_13_n26# ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1651 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1652 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/inv_1/op gnd ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1653 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 ffipg_1/ffi_0/nand_6/a_13_n26# ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1655 gnd ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1656 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a gnd ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1657 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1658 ffipg_1/ffi_0/nand_7/a_13_n26# ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1659 gnd ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1660 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a gnd ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1662 ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1663 ffipg_1/ffi_0/inv_0/op y2in gnd ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1664 ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1665 ffipg_1/ffi_0/inv_1/op clk gnd ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1666 ffipg_1/ffi_1/nand_1/a_13_n26# ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a gnd ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffipg_1/ffi_1/nand_0/a_13_n26# ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 gnd clk ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/inv_0/op gnd ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffipg_1/ffi_1/nand_1/a clk ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 gnd clk ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffipg_1/ffi_1/nand_3/a x2in gnd ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffipg_1/ffi_1/nand_3/a clk ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffipg_1/ffi_1/nand_3/a_13_n26# ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 gnd ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/a gnd ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffipg_1/ffi_1/nand_4/a_13_n26# ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 gnd ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_3/b gnd ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffipg_1/ffi_1/nand_5/a_13_n26# ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/inv_1/op gnd ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffipg_1/ffi_1/nand_6/a_13_n26# ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 gnd ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a gnd ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffipg_1/ffi_1/nand_7/a_13_n26# ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1695 gnd ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1696 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a gnd ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1697 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 ffipg_1/ffi_1/inv_0/op x2in gnd ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 ffipg_1/ffi_1/inv_1/op clk gnd ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 ffipg_2/pggen_0/nand_0/a_13_n26# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1703 gnd ffipg_2/ffi_0/q cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1704 cla_0/l ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1705 cla_0/l ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1706 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1707 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1708 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1709 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 gnd ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1711 ffipg_2/k ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1712 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1713 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1714 ffipg_2/pggen_0/xor_0/a_10_n43# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1715 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1716 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1717 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 cla_2/p0 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1719 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 gnd ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1721 cla_2/p0 ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1722 ffipg_2/ffi_0/nand_1/a_13_n26# ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1723 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1724 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a gnd ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1725 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1726 ffipg_2/ffi_0/nand_0/a_13_n26# ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1727 gnd clk ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1728 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/inv_0/op gnd ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 ffipg_2/ffi_0/nand_1/a clk ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1730 ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1731 gnd clk ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1732 ffipg_2/ffi_0/nand_3/a y3in gnd ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 ffipg_2/ffi_0/nand_3/a clk ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 ffipg_2/ffi_0/nand_3/a_13_n26# ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1735 gnd ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1736 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/a gnd ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1737 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1738 ffipg_2/ffi_0/nand_4/a_13_n26# ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1739 gnd ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1740 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_3/b gnd ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1741 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1742 ffipg_2/ffi_0/nand_5/a_13_n26# ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1743 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1744 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/inv_1/op gnd ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1745 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1746 ffipg_2/ffi_0/nand_6/a_13_n26# ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1747 gnd ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1748 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/a gnd ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1749 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1750 ffipg_2/ffi_0/nand_7/a_13_n26# ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1751 gnd ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1752 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a gnd ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1753 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1754 ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1755 ffipg_2/ffi_0/inv_0/op y3in gnd ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1756 ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1757 ffipg_2/ffi_0/inv_1/op clk gnd ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1758 ffipg_2/ffi_1/nand_1/a_13_n26# ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1759 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1760 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a gnd ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1761 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1762 ffipg_2/ffi_1/nand_0/a_13_n26# ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1763 gnd clk ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1764 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/inv_0/op gnd ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1765 ffipg_2/ffi_1/nand_1/a clk ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1766 ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1767 gnd clk ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1768 ffipg_2/ffi_1/nand_3/a x3in gnd ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1769 ffipg_2/ffi_1/nand_3/a clk ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1770 ffipg_2/ffi_1/nand_3/a_13_n26# ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1771 gnd ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1772 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/a gnd ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1773 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1774 ffipg_2/ffi_1/nand_4/a_13_n26# ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1775 gnd ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1776 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_3/b gnd ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1777 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1778 ffipg_2/ffi_1/nand_5/a_13_n26# ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1779 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1780 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/inv_1/op gnd ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1781 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1782 ffipg_2/ffi_1/nand_6/a_13_n26# ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1783 gnd ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1784 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/a gnd ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1785 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1786 ffipg_2/ffi_1/nand_7/a_13_n26# ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1787 gnd ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1788 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a gnd ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1789 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1790 ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1791 ffipg_2/ffi_1/inv_0/op x3in gnd ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1792 ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1793 ffipg_2/ffi_1/inv_1/op clk gnd ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1794 ffi_1/nand_1/a_13_n26# ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1795 gnd ffi_1/nand_1/b ffi_1/nand_3/b ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1796 ffi_1/nand_3/b ffi_1/nand_1/a gnd ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1797 ffi_1/nand_3/b ffi_1/nand_1/b ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1798 ffi_1/nand_0/a_13_n26# ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1799 gnd clk ffi_1/nand_1/a ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1800 ffi_1/nand_1/a ffi_1/inv_0/op gnd ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1801 ffi_1/nand_1/a clk ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1802 ffi_1/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1803 gnd clk ffi_1/nand_3/a ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1804 ffi_1/nand_3/a cinin gnd ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1805 ffi_1/nand_3/a clk ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1806 ffi_1/nand_3/a_13_n26# ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1807 gnd ffi_1/nand_3/b ffi_1/nand_1/b ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1808 ffi_1/nand_1/b ffi_1/nand_3/a gnd ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1809 ffi_1/nand_1/b ffi_1/nand_3/b ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1810 ffi_1/nand_4/a_13_n26# ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1811 gnd ffi_1/inv_1/op ffi_1/nand_6/a ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1812 ffi_1/nand_6/a ffi_1/nand_3/b gnd ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1813 ffi_1/nand_6/a ffi_1/inv_1/op ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1814 ffi_1/nand_5/a_13_n26# ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1815 gnd ffi_1/nand_1/b ffi_1/nand_7/a ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1816 ffi_1/nand_7/a ffi_1/inv_1/op gnd ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1817 ffi_1/nand_7/a ffi_1/nand_1/b ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1818 ffi_1/nand_6/a_13_n26# ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1819 gnd cinq ffi_1/qbar ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1820 ffi_1/qbar ffi_1/nand_6/a gnd ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1821 ffi_1/qbar cinq ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1822 ffi_1/nand_7/a_13_n26# ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1823 gnd ffi_1/qbar cinq ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1824 cinq ffi_1/nand_7/a gnd ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1825 cinq ffi_1/qbar ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1826 ffi_1/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1827 ffi_1/inv_0/op cinin gnd ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1828 ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1829 ffi_1/inv_1/op clk gnd ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1830 ffi_0/nand_1/a_13_n26# ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1831 gnd ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1832 ffi_0/nand_3/b ffi_0/nand_1/a gnd ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1833 ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1834 ffi_0/nand_0/a_13_n26# ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1835 gnd clk ffi_0/nand_1/a ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1836 ffi_0/nand_1/a ffi_0/inv_0/op gnd ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1837 ffi_0/nand_1/a clk ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1838 ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1839 gnd clk ffi_0/nand_3/a ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1840 ffi_0/nand_3/a cinin gnd ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1841 ffi_0/nand_3/a clk ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1842 ffi_0/nand_3/a_13_n26# ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1843 gnd ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1844 ffi_0/nand_1/b ffi_0/nand_3/a gnd ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1845 ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1846 ffi_0/nand_4/a_13_n26# ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1847 gnd ffi_0/inv_1/op ffi_0/nand_6/a ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1848 ffi_0/nand_6/a ffi_0/nand_3/b gnd ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1849 ffi_0/nand_6/a ffi_0/inv_1/op ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1850 ffi_0/nand_5/a_13_n26# ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1851 gnd ffi_0/nand_1/b ffi_0/nand_7/a ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1852 ffi_0/nand_7/a ffi_0/inv_1/op gnd ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1853 ffi_0/nand_7/a ffi_0/nand_1/b ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1854 ffi_0/nand_6/a_13_n26# ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1855 gnd ffi_0/q nor_0/b ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1856 nor_0/b ffi_0/nand_6/a gnd ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1857 nor_0/b ffi_0/q ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1858 ffi_0/nand_7/a_13_n26# ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1859 gnd nor_0/b ffi_0/q ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1860 ffi_0/q ffi_0/nand_7/a gnd ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1861 ffi_0/q nor_0/b ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1862 ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1863 ffi_0/inv_0/op cinin gnd ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1864 ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1865 ffi_0/inv_1/op clk gnd ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1866 ffipg_3/pggen_0/nand_0/a_13_n26# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1867 gnd ffipg_3/ffi_0/q cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1868 cla_2/g1 ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1869 cla_2/g1 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1870 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1871 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1872 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1873 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1874 gnd ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1875 ffipg_3/k ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1876 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1877 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1878 ffipg_3/pggen_0/xor_0/a_10_n43# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1879 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1880 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1881 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1882 cla_2/p1 ffipg_3/ffi_1/q ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1883 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1884 gnd ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1885 cla_2/p1 ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1886 ffipg_3/ffi_0/nand_1/a_13_n26# ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1887 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1888 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/a gnd ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1889 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1890 ffipg_3/ffi_0/nand_0/a_13_n26# ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1891 gnd clk ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1892 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/inv_0/op gnd ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1893 ffipg_3/ffi_0/nand_1/a clk ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1894 ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1895 gnd clk ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1896 ffipg_3/ffi_0/nand_3/a y4in gnd ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1897 ffipg_3/ffi_0/nand_3/a clk ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1898 ffipg_3/ffi_0/nand_3/a_13_n26# ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1899 gnd ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1900 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/a gnd ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1901 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1902 ffipg_3/ffi_0/nand_4/a_13_n26# ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1903 gnd ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1904 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_3/b gnd ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1905 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1906 ffipg_3/ffi_0/nand_5/a_13_n26# ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1907 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1908 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/inv_1/op gnd ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1909 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1910 ffipg_3/ffi_0/nand_6/a_13_n26# ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1911 gnd ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1912 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/a gnd ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1913 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1914 ffipg_3/ffi_0/nand_7/a_13_n26# ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1915 gnd ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1916 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a gnd ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1917 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1918 ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1919 ffipg_3/ffi_0/inv_0/op y4in gnd ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1920 ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1921 ffipg_3/ffi_0/inv_1/op clk gnd ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1922 ffipg_3/ffi_1/nand_1/a_13_n26# ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1923 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1924 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/a gnd ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1925 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1926 ffipg_3/ffi_1/nand_0/a_13_n26# ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1927 gnd clk ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1928 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/inv_0/op gnd ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1929 ffipg_3/ffi_1/nand_1/a clk ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1930 ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1931 gnd clk ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1932 ffipg_3/ffi_1/nand_3/a x4in gnd ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1933 ffipg_3/ffi_1/nand_3/a clk ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1934 ffipg_3/ffi_1/nand_3/a_13_n26# ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1935 gnd ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1936 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/a gnd ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1937 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1938 ffipg_3/ffi_1/nand_4/a_13_n26# ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1939 gnd ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1940 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_3/b gnd ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1941 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1942 ffipg_3/ffi_1/nand_5/a_13_n26# ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1943 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1944 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/inv_1/op gnd ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1945 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1946 ffipg_3/ffi_1/nand_6/a_13_n26# ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1947 gnd ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1948 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/a gnd ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1949 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1950 ffipg_3/ffi_1/nand_7/a_13_n26# ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1951 gnd ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1952 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a gnd ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1953 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1954 ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1955 ffipg_3/ffi_1/inv_0/op x4in gnd ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1956 ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1957 ffipg_3/ffi_1/inv_1/op clk gnd ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1958 ffipg_5/pggen_0/nand_0/a_13_n26# ffipg_5/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1959 gnd ffipg_5/ffi_0/q ffipg_5/g ffipg_5/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1960 ffipg_5/g ffipg_5/ffi_1/q gnd ffipg_5/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1961 ffipg_5/g ffipg_5/ffi_0/q ffipg_5/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1962 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1963 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/ffi_1/q gnd ffipg_5/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1964 ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1965 ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/ffi_0/q gnd ffipg_5/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1966 gnd ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/a_10_10# ffipg_5/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1967 ffipg_5/k ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1968 gnd ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1969 ffipg_5/pggen_0/xor_0/a_10_10# ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/k ffipg_5/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1970 ffipg_5/pggen_0/xor_0/a_10_n43# ffipg_5/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1971 ffipg_5/pggen_0/xor_0/a_38_n43# ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1972 ffipg_5/pggen_0/xor_0/a_10_10# ffipg_5/ffi_1/q gnd ffipg_5/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1973 ffipg_5/k ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/pggen_0/xor_0/a_10_10# ffipg_5/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1974 ffipg_5/p ffipg_5/ffi_1/q ffipg_5/pggen_0/nor_0/a_13_6# ffipg_5/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1975 ffipg_5/pggen_0/nor_0/a_13_6# ffipg_5/ffi_0/q gnd ffipg_5/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1976 gnd ffipg_5/ffi_1/q ffipg_5/p Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1977 ffipg_5/p ffipg_5/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1978 ffipg_5/ffi_0/nand_1/a_13_n26# ffipg_5/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1979 gnd ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1980 ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_1/a gnd ffipg_5/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1981 ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1982 ffipg_5/ffi_0/nand_0/a_13_n26# ffipg_5/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1983 gnd clk ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1984 ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/inv_0/op gnd ffipg_5/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1985 ffipg_5/ffi_0/nand_1/a clk ffipg_5/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1986 ffipg_5/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1987 gnd clk ffipg_5/ffi_0/nand_3/a ffipg_5/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1988 ffipg_5/ffi_0/nand_3/a y2in gnd ffipg_5/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1989 ffipg_5/ffi_0/nand_3/a clk ffipg_5/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1990 ffipg_5/ffi_0/nand_3/a_13_n26# ffipg_5/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1991 gnd ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1992 ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_3/a gnd ffipg_5/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1993 ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1994 ffipg_5/ffi_0/nand_4/a_13_n26# ffipg_5/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1995 gnd ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_0/nand_6/a ffipg_5/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1996 ffipg_5/ffi_0/nand_6/a ffipg_5/ffi_0/nand_3/b gnd ffipg_5/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1997 ffipg_5/ffi_0/nand_6/a ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1998 ffipg_5/ffi_0/nand_5/a_13_n26# ffipg_5/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1999 gnd ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_7/a ffipg_5/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2000 ffipg_5/ffi_0/nand_7/a ffipg_5/ffi_0/inv_1/op gnd ffipg_5/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2001 ffipg_5/ffi_0/nand_7/a ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2002 ffipg_5/ffi_0/nand_6/a_13_n26# ffipg_5/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2003 gnd ffipg_5/ffi_0/q ffipg_5/ffi_0/qbar ffipg_5/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2004 ffipg_5/ffi_0/qbar ffipg_5/ffi_0/nand_6/a gnd ffipg_5/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2005 ffipg_5/ffi_0/qbar ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2006 ffipg_5/ffi_0/nand_7/a_13_n26# ffipg_5/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2007 gnd ffipg_5/ffi_0/qbar ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2008 ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_7/a gnd ffipg_5/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2009 ffipg_5/ffi_0/q ffipg_5/ffi_0/qbar ffipg_5/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2010 ffipg_5/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2011 ffipg_5/ffi_0/inv_0/op y2in gnd ffipg_5/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2012 ffipg_5/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2013 ffipg_5/ffi_0/inv_1/op clk gnd ffipg_5/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2014 ffipg_5/ffi_1/nand_1/a_13_n26# ffipg_5/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2015 gnd ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2016 ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_1/a gnd ffipg_5/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2017 ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2018 ffipg_5/ffi_1/nand_0/a_13_n26# ffipg_5/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2019 gnd clk ffipg_5/ffi_1/nand_1/a ffipg_5/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2020 ffipg_5/ffi_1/nand_1/a ffipg_5/ffi_1/inv_0/op gnd ffipg_5/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2021 ffipg_5/ffi_1/nand_1/a clk ffipg_5/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2022 ffipg_5/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2023 gnd clk ffipg_5/ffi_1/nand_3/a ffipg_5/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2024 ffipg_5/ffi_1/nand_3/a x2in gnd ffipg_5/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2025 ffipg_5/ffi_1/nand_3/a clk ffipg_5/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2026 ffipg_5/ffi_1/nand_3/a_13_n26# ffipg_5/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2027 gnd ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2028 ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_3/a gnd ffipg_5/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2029 ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2030 ffipg_5/ffi_1/nand_4/a_13_n26# ffipg_5/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2031 gnd ffipg_5/ffi_1/inv_1/op ffipg_5/ffi_1/nand_6/a ffipg_5/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2032 ffipg_5/ffi_1/nand_6/a ffipg_5/ffi_1/nand_3/b gnd ffipg_5/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2033 ffipg_5/ffi_1/nand_6/a ffipg_5/ffi_1/inv_1/op ffipg_5/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2034 ffipg_5/ffi_1/nand_5/a_13_n26# ffipg_5/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2035 gnd ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_7/a ffipg_5/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2036 ffipg_5/ffi_1/nand_7/a ffipg_5/ffi_1/inv_1/op gnd ffipg_5/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2037 ffipg_5/ffi_1/nand_7/a ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2038 ffipg_5/ffi_1/nand_6/a_13_n26# ffipg_5/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2039 gnd ffipg_5/ffi_1/q ffipg_5/ffi_1/qbar ffipg_5/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2040 ffipg_5/ffi_1/qbar ffipg_5/ffi_1/nand_6/a gnd ffipg_5/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2041 ffipg_5/ffi_1/qbar ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2042 ffipg_5/ffi_1/nand_7/a_13_n26# ffipg_5/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2043 gnd ffipg_5/ffi_1/qbar ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2044 ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_7/a gnd ffipg_5/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2045 ffipg_5/ffi_1/q ffipg_5/ffi_1/qbar ffipg_5/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2046 ffipg_5/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2047 ffipg_5/ffi_1/inv_0/op x2in gnd ffipg_5/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2048 ffipg_5/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2049 ffipg_5/ffi_1/inv_1/op clk gnd ffipg_5/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2050 ffipg_4/pggen_0/nand_0/a_13_n26# ffipg_4/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2051 gnd ffipg_4/ffi_0/q ffipg_4/g ffipg_4/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2052 ffipg_4/g ffipg_4/ffi_1/q gnd ffipg_4/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2053 ffipg_4/g ffipg_4/ffi_0/q ffipg_4/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2054 ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2055 ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/ffi_1/q gnd ffipg_4/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2056 ffipg_4/pggen_0/xor_0/inv_1/op ffipg_4/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2057 ffipg_4/pggen_0/xor_0/inv_1/op ffipg_4/ffi_0/q gnd ffipg_4/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2058 gnd ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/a_10_10# ffipg_4/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M2059 ffipg_4/k ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M2060 gnd ffipg_4/pggen_0/xor_0/inv_1/op ffipg_4/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2061 ffipg_4/pggen_0/xor_0/a_10_10# ffipg_4/pggen_0/xor_0/inv_1/op ffipg_4/k ffipg_4/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M2062 ffipg_4/pggen_0/xor_0/a_10_n43# ffipg_4/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2063 ffipg_4/pggen_0/xor_0/a_38_n43# ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2064 ffipg_4/pggen_0/xor_0/a_10_10# ffipg_4/ffi_1/q gnd ffipg_4/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M2065 ffipg_4/k ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/pggen_0/xor_0/a_10_10# ffipg_4/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M2066 p1 ffipg_4/ffi_1/q ffipg_4/pggen_0/nor_0/a_13_6# ffipg_4/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M2067 ffipg_4/pggen_0/nor_0/a_13_6# ffipg_4/ffi_0/q gnd ffipg_4/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M2068 gnd ffipg_4/ffi_1/q p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M2069 p1 ffipg_4/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M2070 ffipg_4/ffi_0/nand_1/a_13_n26# ffipg_4/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2071 gnd ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2072 ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_1/a gnd ffipg_4/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2073 ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2074 ffipg_4/ffi_0/nand_0/a_13_n26# ffipg_4/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2075 gnd clk ffipg_4/ffi_0/nand_1/a ffipg_4/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2076 ffipg_4/ffi_0/nand_1/a ffipg_4/ffi_0/inv_0/op gnd ffipg_4/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2077 ffipg_4/ffi_0/nand_1/a clk ffipg_4/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2078 ffipg_4/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2079 gnd clk ffipg_4/ffi_0/nand_3/a ffipg_4/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2080 ffipg_4/ffi_0/nand_3/a y1in gnd ffipg_4/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2081 ffipg_4/ffi_0/nand_3/a clk ffipg_4/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2082 ffipg_4/ffi_0/nand_3/a_13_n26# ffipg_4/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2083 gnd ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2084 ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_3/a gnd ffipg_4/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2085 ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2086 ffipg_4/ffi_0/nand_4/a_13_n26# ffipg_4/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2087 gnd ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_0/nand_6/a ffipg_4/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2088 ffipg_4/ffi_0/nand_6/a ffipg_4/ffi_0/nand_3/b gnd ffipg_4/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2089 ffipg_4/ffi_0/nand_6/a ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2090 ffipg_4/ffi_0/nand_5/a_13_n26# ffipg_4/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2091 gnd ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_7/a ffipg_4/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2092 ffipg_4/ffi_0/nand_7/a ffipg_4/ffi_0/inv_1/op gnd ffipg_4/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2093 ffipg_4/ffi_0/nand_7/a ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2094 ffipg_4/ffi_0/nand_6/a_13_n26# ffipg_4/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2095 gnd ffipg_4/ffi_0/q ffipg_4/ffi_0/qbar ffipg_4/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2096 ffipg_4/ffi_0/qbar ffipg_4/ffi_0/nand_6/a gnd ffipg_4/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2097 ffipg_4/ffi_0/qbar ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2098 ffipg_4/ffi_0/nand_7/a_13_n26# ffipg_4/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2099 gnd ffipg_4/ffi_0/qbar ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2100 ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_7/a gnd ffipg_4/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2101 ffipg_4/ffi_0/q ffipg_4/ffi_0/qbar ffipg_4/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2102 ffipg_4/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2103 ffipg_4/ffi_0/inv_0/op y1in gnd ffipg_4/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2104 ffipg_4/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2105 ffipg_4/ffi_0/inv_1/op clk gnd ffipg_4/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2106 ffipg_4/ffi_1/nand_1/a_13_n26# ffipg_4/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2107 gnd ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2108 ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_1/a gnd ffipg_4/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2109 ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2110 ffipg_4/ffi_1/nand_0/a_13_n26# ffipg_4/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2111 gnd clk ffipg_4/ffi_1/nand_1/a ffipg_4/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2112 ffipg_4/ffi_1/nand_1/a ffipg_4/ffi_1/inv_0/op gnd ffipg_4/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2113 ffipg_4/ffi_1/nand_1/a clk ffipg_4/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2114 ffipg_4/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2115 gnd clk ffipg_4/ffi_1/nand_3/a ffipg_4/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2116 ffipg_4/ffi_1/nand_3/a x1in gnd ffipg_4/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2117 ffipg_4/ffi_1/nand_3/a clk ffipg_4/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2118 ffipg_4/ffi_1/nand_3/a_13_n26# ffipg_4/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2119 gnd ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2120 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/a gnd ffipg_4/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2121 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2122 ffipg_4/ffi_1/nand_4/a_13_n26# ffipg_4/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2123 gnd ffipg_4/ffi_1/inv_1/op ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2124 ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/nand_3/b gnd ffipg_4/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2125 ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/inv_1/op ffipg_4/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2126 ffipg_4/ffi_1/nand_5/a_13_n26# ffipg_4/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2127 gnd ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2128 ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/inv_1/op gnd ffipg_4/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2129 ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2130 ffipg_4/ffi_1/nand_6/a_13_n26# ffipg_4/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2131 gnd ffipg_4/ffi_1/q ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2132 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_6/a gnd ffipg_4/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2133 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2134 ffipg_4/ffi_1/nand_7/a_13_n26# ffipg_4/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M2135 gnd ffipg_4/ffi_1/qbar ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M2136 ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_7/a gnd ffipg_4/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M2137 ffipg_4/ffi_1/q ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2138 ffipg_4/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2139 ffipg_4/ffi_1/inv_0/op x1in gnd ffipg_4/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M2140 ffipg_4/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M2141 ffipg_4/ffi_1/inv_1/op clk gnd ffipg_4/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 gnd ffipg_2/ffi_0/nand_1/w_0_0# 0.10fF
C1 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C2 gnd ffipg_0/ffi_0/inv_0/op 0.27fF
C3 clk ffo_0/nand_6/a 0.13fF
C4 inv_7/op inv_8/w_0_6# 0.06fF
C5 ffipg_6/ffi_0/nand_1/a ffipg_6/ffi_0/nand_3/b 0.00fF
C6 ffipg_5/p ffipg_5/pggen_0/nand_0/w_0_0# 0.24fF
C7 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar 0.32fF
C8 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/qbar 0.04fF
C9 ffipg_6/ffi_0/nand_6/w_0_0# ffipg_6/ffi_0/nand_6/a 0.06fF
C10 gnd ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C11 x3in ffipg_2/ffi_1/inv_0/op 0.04fF
C12 gnd ffipg_1/ffi_1/nand_1/w_0_0# 0.10fF
C13 clk ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C14 gnd sumffo_3/ffo_0/inv_0/op 0.50fF
C15 sumffo_1/ffo_0/nand_1/b gnd 0.57fF
C16 clk sumffo_0/ffo_0/nand_6/a 0.13fF
C17 cla_2/g1 cla_2/inv_0/in 0.04fF
C18 ffipg_7/ffi_0/nand_2/w_0_0# y4in 0.06fF
C19 ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_0/nand_1/b 0.45fF
C20 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C21 clk ffipg_4/ffi_1/inv_1/op 0.07fF
C22 gnd ffipg_3/ffi_0/nand_7/w_0_0# 0.10fF
C23 gnd nor_1/b 0.34fF
C24 nor_0/w_0_0# inv_0/in 0.11fF
C25 ffipg_7/k ffipg_7/ffi_0/q 0.07fF
C26 ffipg_6/ffi_1/q ffipg_6/pggen_0/xor_0/w_n3_4# 0.06fF
C27 ffi_0/q ffi_0/nand_7/a 0.00fF
C28 ffi_1/inv_1/op cinin 0.01fF
C29 sumffo_1/ffo_0/d sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C30 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C31 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.32fF
C32 gnd ffo_0/d 0.45fF
C33 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C34 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C35 ffipg_6/k gnd 0.27fF
C36 ffipg_5/ffi_0/q ffipg_5/pggen_0/nand_0/w_0_0# 0.06fF
C37 ffipg_3/ffi_1/nand_2/w_0_0# ffipg_3/ffi_1/nand_3/a 0.04fF
C38 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_3/b 0.00fF
C39 ffipg_7/ffi_1/nand_7/w_0_0# ffipg_7/ffi_1/nand_7/a 0.06fF
C40 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_3/b 0.04fF
C41 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C42 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/pggen_0/xor_0/inv_1/op 0.08fF
C43 cla_1/l cla_0/n 0.01fF
C44 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a 0.31fF
C45 nor_4/a nor_4/w_0_0# 0.07fF
C46 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C47 ffipg_6/ffi_0/qbar ffipg_6/ffi_0/nand_7/w_0_0# 0.06fF
C48 ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_6/w_0_0# 0.06fF
C49 gnd ffipg_4/ffi_0/nand_1/a 0.44fF
C50 gnd ffipg_3/ffi_1/nand_4/w_0_0# 0.10fF
C51 gnd ffipg_2/ffi_1/nand_7/w_0_0# 0.10fF
C52 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a 0.31fF
C53 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/a 0.06fF
C54 gnd ffipg_1/ffi_0/inv_0/op 0.27fF
C55 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_5/w_0_0# 0.06fF
C56 ffipg_6/ffi_1/q ffipg_6/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C57 y4in ffipg_3/ffi_0/inv_1/op 0.01fF
C58 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C59 gnd ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C60 gnd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C61 ffipg_7/ffi_1/inv_0/op x4in 0.04fF
C62 ffipg_7/pggen_0/xor_0/inv_0/op gnd 0.32fF
C63 ffipg_5/ffi_1/q ffipg_5/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C64 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_3/b 0.04fF
C65 ffi_1/qbar ffi_1/nand_7/a 0.31fF
C66 ffi_1/nand_6/a cinq 0.31fF
C67 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/inv_1/w_0_6# 0.04fF
C68 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a 0.31fF
C69 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C70 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_1/b 0.04fF
C71 gnd sumffo_3/ffo_0/nand_1/a 0.33fF
C72 gnd sumffo_2/ffo_0/nand_1/w_0_0# 0.10fF
C73 ffipg_4/ffi_1/inv_0/op ffipg_4/ffi_1/nand_0/w_0_0# 0.06fF
C74 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_6/a 0.04fF
C75 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C76 clk ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C77 ffo_0/inv_0/op ffo_0/inv_0/w_0_6# 0.03fF
C78 ffipg_7/ffi_1/inv_1/w_0_6# clk 0.06fF
C79 ffipg_6/ffi_0/nand_2/w_0_0# clk 0.06fF
C80 ffipg_4/ffi_0/q ffipg_4/k 0.07fF
C81 gnd ffipg_4/ffi_0/nand_7/w_0_0# 0.10fF
C82 ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/nand_0/w_0_0# 0.04fF
C83 clk ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C84 inv_0/in nor_0/b 0.16fF
C85 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C86 sumffo_0/ffo_0/nand_0/a_13_n26# gnd 0.01fF
C87 ffipg_7/pggen_0/xor_0/w_n3_4# ffipg_7/ffi_0/q 0.06fF
C88 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C89 gnd ffipg_1/ffi_1/inv_1/op 1.85fF
C90 gnd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C91 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C92 gnd ffipg_3/k 0.61fF
C93 ffipg_7/pggen_0/nand_0/w_0_0# ffipg_7/ffi_1/q 0.06fF
C94 ffipg_7/ffi_0/qbar ffipg_7/ffi_0/nand_7/w_0_0# 0.06fF
C95 ffipg_0/k nor_0/b 0.06fF
C96 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/inv_1/w_0_6# 0.04fF
C97 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C98 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C99 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C100 clk ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C101 gnd ffipg_1/ffi_1/nand_7/a 0.37fF
C102 gnd inv_7/in 0.43fF
C103 gnd inv_2/in 0.47fF
C104 ffipg_7/ffi_1/nand_4/w_0_0# ffipg_7/ffi_1/nand_3/b 0.06fF
C105 ffipg_6/g gnd 0.31fF
C106 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C107 gnd ffipg_5/ffi_0/inv_1/w_0_6# 0.06fF
C108 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/qbar 0.00fF
C109 gnd ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C110 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C111 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a 0.13fF
C112 gnd sumffo_3/ffo_0/nand_2/w_0_0# 0.10fF
C113 inv_7/op ffi_0/q 0.31fF
C114 ffipg_7/ffi_1/nand_6/a ffipg_7/ffi_1/qbar 0.00fF
C115 ffipg_7/g ffipg_7/ffi_0/q 0.13fF
C116 x3in ffipg_2/ffi_1/inv_1/op 0.01fF
C117 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/a 0.06fF
C118 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# 0.04fF
C119 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/b 0.31fF
C120 gnd ffipg_4/ffi_1/nand_7/a 0.37fF
C121 clk ffipg_5/ffi_0/inv_0/op 0.32fF
C122 y3in ffipg_2/ffi_0/inv_0/op 0.04fF
C123 gnd ffipg_2/ffi_0/nand_2/w_0_0# 0.10fF
C124 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/ffi_1/q 0.06fF
C125 gnd sumffo_2/ffo_0/nand_5/w_0_0# 0.10fF
C126 ffipg_7/pggen_0/xor_0/inv_1/op gnd 0.35fF
C127 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/inv_0/op 0.06fF
C128 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C129 cla_0/inv_0/in cla_0/l 0.07fF
C130 ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_7/a 0.00fF
C131 clk ffipg_4/ffi_0/inv_0/op 0.32fF
C132 gnd ffipg_5/ffi_1/inv_1/w_0_6# 0.06fF
C133 ffipg_5/ffi_0/nand_1/w_0_0# ffipg_5/ffi_0/nand_1/b 0.06fF
C134 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/nand_7/a 0.06fF
C135 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/inv_1/op 0.33fF
C136 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C137 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_3/b 0.00fF
C138 ffipg_4/pggen_0/nor_0/w_0_0# ffipg_4/k 0.21fF
C139 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C140 gnd nor_3/b 0.33fF
C141 ffi_0/q inv_8/w_0_6# 0.06fF
C142 ffipg_7/k ffipg_7/p 0.05fF
C143 ffipg_6/ffi_1/nand_3/b gnd 0.74fF
C144 gnd ffipg_5/ffi_1/nand_3/w_0_0# 0.11fF
C145 gnd ffi_0/nand_1/a 0.44fF
C146 ffi_1/nand_3/w_0_0# ffi_1/nand_3/a 0.06fF
C147 clk ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C148 ffipg_2/ffi_0/inv_0/op ffipg_2/ffi_0/inv_0/w_0_6# 0.03fF
C149 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_0/q 0.12fF
C150 cla_0/g0 ffipg_0/ffi_0/q 0.13fF
C151 clk sumffo_1/ffo_0/nand_0/b 0.04fF
C152 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C153 cla_2/l cla_2/p1 0.02fF
C154 ffipg_7/ffi_1/nand_1/w_0_0# gnd 0.10fF
C155 ffipg_6/ffi_0/nand_4/w_0_0# ffipg_6/ffi_0/inv_1/op 0.06fF
C156 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a 0.31fF
C157 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_1/b 0.04fF
C158 clk ffo_0/inv_1/w_0_6# 0.06fF
C159 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/inv_1/op 0.33fF
C160 gnd p1 0.35fF
C161 clk ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C162 gnd ffipg_3/ffi_1/nand_6/a 0.37fF
C163 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/qbar 0.00fF
C164 gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C165 ffi_1/inv_0/op cinin 0.04fF
C166 ffo_0/d ffo_0/nand_0/b 0.40fF
C167 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C168 sumffo_1/ffo_0/nand_6/a sumffo_1/sbar 0.00fF
C169 cla_0/g0 cla_0/inv_0/in 0.16fF
C170 x4in ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C171 ffipg_6/ffi_1/inv_1/w_0_6# clk 0.06fF
C172 ffipg_3/ffi_0/inv_0/op y4in 0.04fF
C173 ffi_0/q sumffo_2/ffo_0/d 0.27fF
C174 clk ffipg_5/ffi_1/nand_0/w_0_0# 0.06fF
C175 gnd ffipg_5/ffi_0/nand_6/w_0_0# 0.10fF
C176 gnd ffipg_1/ffi_1/nand_3/b 0.74fF
C177 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/ffi_0/q 0.06fF
C178 gnd ffipg_0/ffi_1/nand_1/a 0.44fF
C179 inv_1/in nor_1/w_0_0# 0.11fF
C180 ffo_0/nand_6/w_0_0# ffo_0/qbar 0.04fF
C181 ffo_0/nand_1/b ffo_0/nand_7/a 0.13fF
C182 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C183 sumffo_0/sbar z1o 0.32fF
C184 ffipg_7/ffi_0/nand_5/w_0_0# ffipg_7/ffi_0/nand_7/a 0.04fF
C185 ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/nand_4/w_0_0# 0.06fF
C186 ffipg_4/ffi_1/q ffipg_4/pggen_0/xor_0/w_n3_4# 0.06fF
C187 ffipg_5/ffi_1/nand_1/w_0_0# ffipg_5/ffi_1/nand_1/a 0.06fF
C188 ffipg_6/ffi_1/nand_2/w_0_0# gnd 0.10fF
C189 ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_6/a 0.31fF
C190 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/a 0.06fF
C191 sumffo_1/ffo_0/nand_6/a z2o 0.31fF
C192 cla_2/inv_0/w_0_6# gnd 0.06fF
C193 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C194 ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/k 0.52fF
C195 gnd ffipg_5/ffi_1/nand_6/w_0_0# 0.10fF
C196 ffipg_5/ffi_0/nand_4/w_0_0# ffipg_5/ffi_0/nand_3/b 0.06fF
C197 ffi_0/nand_7/w_0_0# ffi_0/nand_7/a 0.06fF
C198 gnd ffipg_2/ffi_1/nand_4/w_0_0# 0.10fF
C199 gnd ffipg_1/ffi_1/nand_0/w_0_0# 0.10fF
C200 ffipg_0/ffi_0/q ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C201 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C202 nand_2/b inv_3/w_0_6# 0.06fF
C203 gnd ffipg_2/ffi_0/nand_1/a 0.44fF
C204 gnd ffo_0/nand_5/w_0_0# 0.10fF
C205 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C206 ffipg_2/ffi_1/nand_7/w_0_0# ffipg_2/ffi_1/nand_7/a 0.06fF
C207 ffipg_5/ffi_1/nand_1/a ffipg_5/ffi_1/nand_3/b 0.00fF
C208 clk ffipg_4/ffi_1/nand_1/a 0.13fF
C209 gnd ffipg_5/ffi_1/nand_3/a 0.33fF
C210 clk ffipg_3/ffi_0/nand_1/a 0.13fF
C211 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.35fF
C212 ffipg_0/ffi_0/nand_2/w_0_0# ffipg_0/ffi_0/nand_3/a 0.04fF
C213 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C214 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C215 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C216 sumffo_0/ffo_0/nand_5/w_0_0# gnd 0.10fF
C217 ffipg_6/ffi_0/nand_3/w_0_0# gnd 0.11fF
C218 ffipg_4/ffi_0/nand_2/w_0_0# ffipg_4/ffi_0/nand_3/a 0.04fF
C219 ffipg_5/ffi_1/nand_3/a ffipg_5/ffi_1/nand_3/w_0_0# 0.06fF
C220 ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_1/inv_1/op 0.75fF
C221 gnd ffipg_2/ffi_1/nand_0/a_13_n26# 0.01fF
C222 ffi_0/q sumffo_1/xor_0/inv_1/op 0.04fF
C223 ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_7/w_0_0# 0.04fF
C224 gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C225 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C226 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op 0.06fF
C227 y4in ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C228 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/inv_1/op 0.06fF
C229 gnd ffipg_0/ffi_1/inv_0/op 0.27fF
C230 ffipg_0/pggen_0/nand_0/w_0_0# ffipg_0/ffi_1/q 0.06fF
C231 clk ffipg_0/ffi_0/nand_1/a 0.13fF
C232 cla_0/g0 nor_0/w_0_0# 0.06fF
C233 ffipg_7/ffi_1/nand_3/a gnd 0.33fF
C234 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_1/b 0.04fF
C235 ffi_1/nand_1/b ffi_1/nand_1/w_0_0# 0.06fF
C236 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/qbar 0.00fF
C237 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_3/b 0.00fF
C238 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C239 gnd ffi_1/nand_5/w_0_0# 0.10fF
C240 gnd ffipg_1/ffi_1/nand_1/a 0.44fF
C241 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C242 gnd sumffo_1/ffo_0/nand_3/w_0_0# 0.11fF
C243 sumffo_0/xor_0/inv_1/op gnd 0.35fF
C244 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C245 ffipg_6/ffi_1/nand_0/w_0_0# clk 0.06fF
C246 ffipg_5/ffi_1/inv_1/op ffipg_5/ffi_1/inv_1/w_0_6# 0.04fF
C247 gnd ffipg_3/ffi_0/nand_7/a 0.37fF
C248 ffipg_7/ffi_1/nand_2/w_0_0# gnd 0.10fF
C249 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C250 ffipg_4/ffi_1/nand_3/b ffipg_4/ffi_1/inv_1/op 0.33fF
C251 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_1/a 0.06fF
C252 nor_3/w_0_0# cla_2/n 0.06fF
C253 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C254 gnd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C255 cla_0/l cla_2/g1 0.26fF
C256 cla_1/nand_0/w_0_0# gnd 0.10fF
C257 ffipg_7/ffi_1/nand_1/w_0_0# ffipg_7/ffi_1/nand_3/b 0.04fF
C258 ffipg_7/ffi_1/nand_3/b gnd 0.74fF
C259 ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/w_n3_4# 0.06fF
C260 gnd ffipg_5/ffi_1/inv_1/op 1.85fF
C261 gnd ffipg_5/ffi_0/nand_3/w_0_0# 0.11fF
C262 gnd ffi_0/nand_3/w_0_0# 0.11fF
C263 gnd ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C264 inv_8/w_0_6# inv_8/in 0.10fF
C265 gnd ffo_0/nand_0/b 0.58fF
C266 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d 0.04fF
C267 cla_2/g1 cla_2/n 0.13fF
C268 ffipg_7/pggen_0/xor_0/a_10_10# gnd 0.93fF
C269 ffipg_6/ffi_0/nand_0/w_0_0# clk 0.06fF
C270 cla_0/n inv_3/w_0_6# 0.14fF
C271 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C272 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C273 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/xor_0/inv_0/op 0.03fF
C274 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C275 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C276 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C277 ffipg_4/ffi_0/nand_4/w_0_0# ffipg_4/ffi_0/inv_1/op 0.06fF
C278 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_3/b 0.00fF
C279 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a 0.31fF
C280 nor_4/a inv_9/in 0.02fF
C281 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C282 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C283 ffi_0/q ffipg_1/k 0.06fF
C284 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_7/w_0_0# 0.06fF
C285 gnd ffipg_5/g 0.31fF
C286 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C287 gnd sumffo_2/ffo_0/inv_0/w_0_6# 0.07fF
C288 sumffo_0/xor_0/w_n3_4# gnd 0.12fF
C289 ffipg_7/ffi_1/inv_0/w_0_6# gnd 0.06fF
C290 ffipg_4/ffi_1/nand_3/w_0_0# ffipg_4/ffi_1/nand_3/a 0.06fF
C291 gnd ffipg_4/pggen_0/xor_0/inv_1/op 0.35fF
C292 gnd ffipg_5/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C293 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C294 gnd ffipg_2/ffi_1/nand_7/a 0.37fF
C295 gnd ffipg_2/ffi_0/q 3.00fF
C296 gnd ffipg_1/ffi_1/nand_6/w_0_0# 0.10fF
C297 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/b 0.31fF
C298 clk ffi_1/nand_2/w_0_0# 0.06fF
C299 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_0/w_0_0# 0.04fF
C300 clk ffipg_0/ffi_0/inv_0/op 0.32fF
C301 gnd ffipg_0/ffi_1/q 2.24fF
C302 ffipg_6/pggen_0/xor_0/inv_1/op gnd 0.35fF
C303 ffipg_5/ffi_1/q ffipg_5/ffi_1/qbar 0.32fF
C304 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C305 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/w_0_0# 0.06fF
C306 gnd ffipg_4/ffi_0/nand_5/w_0_0# 0.10fF
C307 ffipg_1/ffi_0/nand_7/w_0_0# ffipg_1/ffi_0/nand_7/a 0.06fF
C308 gnd ffipg_0/ffi_0/nand_5/w_0_0# 0.10fF
C309 gnd sumffo_3/ffo_0/nand_3/b 0.74fF
C310 cla_1/inv_0/in gnd 0.34fF
C311 ffipg_7/ffi_1/qbar ffipg_7/ffi_1/nand_7/w_0_0# 0.06fF
C312 ffipg_7/ffi_0/q ffipg_7/p 0.03fF
C313 ffipg_6/ffi_0/nand_6/a gnd 0.37fF
C314 sumffo_1/ffo_0/nand_1/b clk 0.45fF
C315 ffipg_6/ffi_0/nand_2/w_0_0# ffipg_6/ffi_0/nand_3/a 0.04fF
C316 gnd ffipg_2/ffi_0/nand_5/w_0_0# 0.10fF
C317 ffipg_2/k ffipg_2/ffi_1/q 0.46fF
C318 gnd ffipg_0/ffi_0/nand_7/w_0_0# 0.10fF
C319 gnd sumffo_2/sbar 0.62fF
C320 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_6/a 0.04fF
C321 cla_0/inv_0/in cla_1/p0 0.02fF
C322 ffipg_7/ffi_1/nand_7/a gnd 0.37fF
C323 gnd ffi_1/nand_0/w_0_0# 0.10fF
C324 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C325 ffipg_4/ffi_0/nand_6/w_0_0# ffipg_4/ffi_0/qbar 0.04fF
C326 ffipg_5/k ffipg_5/pggen_0/xor_0/a_10_10# 0.45fF
C327 ffipg_0/ffi_1/nand_4/w_0_0# ffipg_0/ffi_1/nand_6/a 0.04fF
C328 inv_0/op nor_0/w_0_0# 0.10fF
C329 gnd ffi_1/nand_7/w_0_0# 0.10fF
C330 gnd ffipg_1/ffi_0/nand_7/a 0.37fF
C331 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_1/b 0.06fF
C332 ffipg_0/ffi_1/nand_6/w_0_0# ffipg_0/ffi_1/qbar 0.04fF
C333 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_3/b 0.04fF
C334 gnd ffipg_0/ffi_0/nand_3/b 0.74fF
C335 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_3/a 0.04fF
C336 gnd sumffo_2/ffo_0/inv_0/op 0.50fF
C337 ffipg_7/ffi_1/nand_2/w_0_0# ffipg_7/ffi_1/nand_3/a 0.04fF
C338 ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_0/inv_1/w_0_6# 0.04fF
C339 ffipg_6/ffi_1/nand_7/w_0_0# ffipg_6/ffi_1/nand_7/a 0.06fF
C340 ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_1/inv_1/op 0.75fF
C341 ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/k 0.52fF
C342 gnd ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C343 gnd couto 0.80fF
C344 ffipg_7/ffi_1/nand_3/a ffipg_7/ffi_1/nand_3/b 0.31fF
C345 sumffo_0/ffo_0/inv_0/op gnd 0.27fF
C346 ffipg_7/ffi_0/nand_1/a ffipg_7/ffi_0/nand_1/b 0.31fF
C347 ffipg_6/ffi_1/nand_5/w_0_0# ffipg_6/ffi_1/nand_7/a 0.04fF
C348 clk ffipg_4/ffi_0/nand_1/a 0.13fF
C349 clk ffipg_1/ffi_0/inv_0/op 0.32fF
C350 ffipg_7/pggen_0/nand_0/w_0_0# ffipg_7/g 0.04fF
C351 ffo_0/qbar ffo_0/nand_7/a 0.31fF
C352 gnd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C353 ffi_0/q inv_8/in 0.13fF
C354 ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_6/w_0_0# 0.06fF
C355 gnd ffipg_5/ffi_1/nand_0/a_13_n26# 0.01fF
C356 x2in ffipg_5/ffi_1/inv_0/w_0_6# 0.06fF
C357 ffipg_3/ffi_1/inv_0/op ffipg_3/ffi_1/inv_0/w_0_6# 0.03fF
C358 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a 0.13fF
C359 gnd sumffo_3/ffo_0/nand_3/a 0.33fF
C360 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C361 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a 0.13fF
C362 ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_7/w_0_0# 0.04fF
C363 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C364 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C365 sumffo_3/ffo_0/d sumffo_3/ffo_0/inv_0/w_0_6# 0.06fF
C366 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C367 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C368 gnd ffi_0/inv_1/w_0_6# 0.06fF
C369 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/qbar 0.04fF
C370 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a 0.13fF
C371 clk ffipg_1/ffi_1/inv_1/op 0.07fF
C372 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C373 gnd ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C374 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# 0.04fF
C375 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/k 0.06fF
C376 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/inv_1/op 0.33fF
C377 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_1/b 0.31fF
C378 ffi_0/q sumffo_1/xor_0/w_n3_4# 0.00fF
C379 clk ffipg_5/ffi_0/inv_1/w_0_6# 0.06fF
C380 gnd ffipg_5/ffi_0/nand_6/a 0.37fF
C381 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/qbar 0.04fF
C382 ffi_0/q ffi_0/nand_7/w_0_0# 0.04fF
C383 ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# 0.04fF
C384 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C385 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/nand_6/a 0.04fF
C386 inv_0/in nor_0/a 0.02fF
C387 ffo_0/nand_6/a ffo_0/qbar 0.00fF
C388 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C389 sumffo_0/sbar gnd 0.62fF
C390 cla_0/l cla_1/inv_0/op 0.35fF
C391 ffipg_7/ffi_1/nand_0/w_0_0# gnd 0.10fF
C392 clk ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C393 ffipg_0/k nor_0/a 0.05fF
C394 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C395 clk sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C396 gnd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C397 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_5/w_0_0# 0.06fF
C398 ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C399 clk ffipg_5/ffi_1/inv_1/w_0_6# 0.06fF
C400 gnd ffipg_5/ffi_1/nand_6/a 0.37fF
C401 ffipg_5/pggen_0/nor_0/w_0_0# ffipg_5/p 0.05fF
C402 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C403 ffi_0/nand_1/a ffi_0/nand_3/b 0.00fF
C404 gnd ffi_0/nand_3/b 0.74fF
C405 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C406 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C407 gnd ffipg_2/ffi_0/nand_3/a 0.33fF
C408 ffipg_4/ffi_0/inv_0/op ffipg_4/ffi_0/inv_0/w_0_6# 0.03fF
C409 y2in ffipg_5/ffi_0/inv_0/op 0.04fF
C410 ffipg_7/pggen_0/nand_0/w_0_0# ffipg_7/ffi_0/q 0.06fF
C411 ffipg_4/ffi_0/inv_0/op ffipg_4/ffi_0/nand_0/w_0_0# 0.06fF
C412 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_6/w_0_0# 0.04fF
C413 gnd ffipg_4/ffi_0/nand_0/a_13_n26# 0.01fF
C414 gnd ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C415 gnd ffipg_4/ffi_0/q 3.00fF
C416 ffipg_5/ffi_0/nand_6/w_0_0# ffipg_5/ffi_0/nand_6/a 0.06fF
C417 clk ffi_0/nand_1/a 0.13fF
C418 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C419 ffipg_7/ffi_1/nand_5/w_0_0# ffipg_7/ffi_1/nand_1/b 0.06fF
C420 ffipg_7/ffi_0/inv_1/op y4in 0.01fF
C421 clk gnd 34.68fF
C422 ffipg_4/ffi_1/nand_1/a ffipg_4/ffi_1/nand_3/b 0.00fF
C423 gnd ffipg_4/ffi_1/nand_3/a 0.33fF
C424 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C425 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C426 gnd sumffo_3/ffo_0/nand_6/a 0.33fF
C427 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C428 sumffo_2/ffo_0/nand_7/w_0_0# z3o 0.04fF
C429 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C430 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_4/w_0_0# 0.06fF
C431 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/inv_1/op 0.45fF
C432 ffipg_6/ffi_1/nand_1/w_0_0# ffipg_6/ffi_1/nand_3/b 0.04fF
C433 gnd ffi_0/nand_0/a_13_n26# 0.01fF
C434 ffipg_4/ffi_0/q p1 0.03fF
C435 ffipg_5/ffi_1/nand_0/w_0_0# ffipg_5/ffi_1/inv_0/op 0.06fF
C436 ffipg_5/pggen_0/nor_0/w_0_0# ffipg_5/ffi_0/q 0.06fF
C437 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C438 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/nand_6/a 0.04fF
C439 ffi_1/nand_3/w_0_0# ffi_1/nand_3/b 0.06fF
C440 ffipg_1/ffi_1/nand_2/w_0_0# x2in 0.06fF
C441 ffipg_0/pggen_0/nand_0/w_0_0# ffipg_0/ffi_0/q 0.06fF
C442 gnd ffipg_2/ffi_0/nand_0/a_13_n26# 0.01fF
C443 ffipg_1/k ffipg_1/ffi_0/q 0.07fF
C444 gnd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C445 ffipg_6/ffi_1/nand_1/w_0_0# gnd 0.10fF
C446 ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_6/a 0.31fF
C447 ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/k 0.06fF
C448 ffipg_5/ffi_1/nand_6/w_0_0# ffipg_5/ffi_1/nand_6/a 0.06fF
C449 gnd ffipg_5/pggen_0/xor_0/a_10_10# 0.93fF
C450 cinin ffi_0/inv_0/w_0_6# 0.06fF
C451 ffi_0/q ffi_0/nand_6/w_0_0# 0.06fF
C452 ffi_1/inv_1/op ffi_1/nand_3/b 0.33fF
C453 clk ffipg_0/ffi_1/nand_1/a 0.13fF
C454 gnd sumffo_1/ffo_0/nand_3/a 0.48fF
C455 ffipg_7/ffi_0/nand_0/w_0_0# gnd 0.10fF
C456 ffipg_6/ffi_0/inv_0/op ffipg_6/ffi_0/inv_0/w_0_6# 0.03fF
C457 ffipg_6/ffi_1/nand_2/w_0_0# clk 0.06fF
C458 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C459 gnd ffipg_4/ffi_0/inv_1/w_0_6# 0.06fF
C460 ffo_0/d nor_4/w_0_0# 0.03fF
C461 gnd ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C462 sumffo_1/sbar sumffo_1/ffo_0/nand_7/w_0_0# 0.06fF
C463 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C464 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/inv_0/w_0_6# 0.03fF
C465 inv_6/in cla_2/n 0.02fF
C466 gnd sumffo_3/ffo_0/nand_6/w_0_0# 0.10fF
C467 ffipg_4/ffi_0/nand_7/w_0_0# ffipg_4/ffi_0/nand_7/a 0.06fF
C468 gnd ffipg_4/pggen_0/nor_0/w_0_0# 0.11fF
C469 gnd ffipg_5/pggen_0/xor_0/inv_1/op 0.35fF
C470 gnd ffi_0/nand_3/a 0.33fF
C471 clk ffipg_1/ffi_1/nand_0/w_0_0# 0.06fF
C472 clk ffipg_2/ffi_0/nand_1/a 0.13fF
C473 clk ffo_0/nand_5/w_0_0# 0.06fF
C474 ffipg_5/ffi_1/nand_0/w_0_0# ffipg_5/ffi_1/nand_1/a 0.04fF
C475 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C476 ffi_1/inv_0/op ffi_1/inv_0/w_0_6# 0.03fF
C477 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_1/b 0.45fF
C478 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C479 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b 0.13fF
C480 ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/inv_1/op 0.33fF
C481 ffipg_4/pggen_0/nor_0/w_0_0# p1 0.05fF
C482 clk ffipg_5/ffi_1/nand_3/a 0.13fF
C483 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C484 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_1/b 0.04fF
C485 ffi_0/nand_2/w_0_0# cinin 0.06fF
C486 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C487 sumffo_0/ffo_0/nand_5/w_0_0# clk 0.06fF
C488 ffipg_7/ffi_0/inv_0/op gnd 0.27fF
C489 ffipg_6/ffi_0/qbar ffipg_6/ffi_0/nand_7/a 0.31fF
C490 ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_0/nand_6/a 0.13fF
C491 ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C492 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a 0.13fF
C493 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a 0.13fF
C494 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C495 gnd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C496 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/d 0.40fF
C497 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/nand_3/a 0.04fF
C498 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C499 ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_6/a 0.31fF
C500 ffipg_4/ffi_1/nand_3/w_0_0# ffipg_4/ffi_1/nand_3/b 0.06fF
C501 ffi_0/q sumffo_3/xor_0/w_n3_4# 0.01fF
C502 clk ffipg_0/ffi_1/inv_0/op 0.32fF
C503 nor_2/w_0_0# nor_2/b 0.06fF
C504 ffipg_6/ffi_1/q ffipg_6/pggen_0/nor_0/w_0_0# 0.06fF
C505 ffi_0/inv_0/op ffi_0/inv_0/w_0_6# 0.03fF
C506 ffi_0/q ffi_0/nand_6/a 0.31fF
C507 nor_4/b nor_4/a 0.42fF
C508 gnd ffipg_0/ffi_0/q 3.00fF
C509 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C510 inv_1/op ffipg_2/k 0.09fF
C511 cla_2/nor_0/w_0_0# cla_2/p0 0.06fF
C512 cla_0/l inv_2/w_0_6# 0.06fF
C513 ffipg_7/ffi_1/nand_3/a clk 0.13fF
C514 ffipg_7/ffi_0/nand_1/a gnd 0.44fF
C515 gnd ffipg_4/g 0.31fF
C516 gnd ffi_0/nand_5/w_0_0# 0.10fF
C517 gnd ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C518 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op 0.06fF
C519 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/b 0.31fF
C520 gnd sumffo_2/xor_0/inv_0/op 0.32fF
C521 inv_3/in inv_3/w_0_6# 0.10fF
C522 ffipg_6/ffi_1/nand_7/w_0_0# gnd 0.10fF
C523 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_6/a 0.00fF
C524 ffipg_5/ffi_1/inv_1/op ffipg_5/ffi_1/nand_6/a 0.13fF
C525 ffi_0/inv_1/op cinin 0.01fF
C526 ffi_0/nand_3/w_0_0# ffi_0/nand_3/b 0.06fF
C527 clk ffipg_1/ffi_1/nand_1/a 0.13fF
C528 ffipg_7/ffi_1/nand_2/w_0_0# clk 0.06fF
C529 ffipg_6/ffi_1/nand_5/w_0_0# gnd 0.10fF
C530 cla_2/l inv_5/in 0.05fF
C531 gnd ffipg_4/ffi_0/nand_7/a 0.37fF
C532 gnd ffipg_5/pggen_0/xor_0/inv_0/op 0.32fF
C533 gnd ffipg_2/ffi_0/inv_1/op 1.85fF
C534 gnd ffipg_0/ffi_0/nand_7/a 0.37fF
C535 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a 0.31fF
C536 gnd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C537 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a 0.31fF
C538 ffipg_6/ffi_0/inv_0/op y3in 0.04fF
C539 gnd ffipg_1/ffi_1/nand_1/b 0.57fF
C540 cla_0/inv_0/in gnd 0.34fF
C541 ffipg_7/pggen_0/nand_0/w_0_0# ffipg_7/p 0.24fF
C542 gnd ffipg_5/ffi_0/nand_4/w_0_0# 0.10fF
C543 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C544 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.35fF
C545 ffipg_3/pggen_0/nand_0/w_0_0# ffipg_3/ffi_0/q 0.06fF
C546 cla_1/inv_0/w_0_6# cla_0/n 0.23fF
C547 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C548 ffipg_7/ffi_0/qbar ffipg_7/ffi_0/nand_7/a 0.31fF
C549 clk ffipg_5/ffi_1/inv_1/op 0.07fF
C550 ffipg_5/k ffipg_5/pggen_0/nor_0/a_13_6# 0.01fF
C551 clk ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C552 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a 0.31fF
C553 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/qbar 0.04fF
C554 inv_1/op nor_1/w_0_0# 0.03fF
C555 clk ffo_0/nand_0/b 0.04fF
C556 gnd sumffo_3/xor_0/inv_1/op 0.35fF
C557 cla_1/l inv_3/w_0_6# 0.06fF
C558 ffipg_3/ffi_1/q ffipg_3/ffi_0/q 0.73fF
C559 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C560 ffi_1/nand_6/w_0_0# ffi_1/qbar 0.04fF
C561 gnd ffi_1/nand_7/a 0.33fF
C562 gnd ffipg_1/ffi_1/nand_3/w_0_0# 0.11fF
C563 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/qbar 0.00fF
C564 gnd ffipg_0/ffi_1/nand_3/b 0.74fF
C565 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/a 0.06fF
C566 ffi_0/inv_1/op ffi_0/nand_6/a 0.13fF
C567 ffi_0/inv_0/op ffi_0/nand_0/w_0_0# 0.06fF
C568 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C569 ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/nand_3/b 0.00fF
C570 gnd ffipg_3/ffi_0/nand_3/a 0.33fF
C571 gnd ffipg_2/ffi_1/nand_5/w_0_0# 0.10fF
C572 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/ffi_1/q 0.06fF
C573 gnd ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C574 gnd sumffo_2/ffo_0/nand_1/b 0.57fF
C575 cla_0/l nor_0/a 0.16fF
C576 gnd nor_4/w_0_0# 0.15fF
C577 ffo_0/nand_3/w_0_0# ffo_0/nand_3/a 0.06fF
C578 sumffo_0/ffo_0/nand_1/a gnd 0.44fF
C579 cla_2/l cla_0/l 0.37fF
C580 ffipg_7/ffi_1/qbar gnd 0.67fF
C581 ffipg_6/ffi_1/nand_4/w_0_0# ffipg_6/ffi_1/inv_1/op 0.06fF
C582 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/inv_1/op 0.45fF
C583 ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/inv_1/op 0.22fF
C584 gnd ffi_0/nand_1/w_0_0# 0.10fF
C585 ffi_0/nand_1/w_0_0# ffi_0/nand_1/a 0.06fF
C586 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b 0.32fF
C587 ffipg_6/ffi_0/nand_7/w_0_0# ffipg_6/ffi_0/nand_7/a 0.06fF
C588 gnd ffipg_1/ffi_1/qbar 0.67fF
C589 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_1/inv_1/op 0.75fF
C590 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar 0.32fF
C591 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C592 gnd ffipg_1/ffi_0/nand_6/w_0_0# 0.10fF
C593 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_3/b 0.00fF
C594 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C595 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C596 gnd sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C597 ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/inv_1/op 0.33fF
C598 ffipg_7/ffi_1/q ffipg_7/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C599 inv_1/op inv_1/in 0.04fF
C600 ffi_0/nand_3/w_0_0# ffi_0/nand_3/a 0.06fF
C601 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C602 cla_0/l nand_2/b 0.06fF
C603 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C604 cla_0/g0 nor_0/a 0.68fF
C605 clk ffi_1/nand_0/w_0_0# 0.06fF
C606 gnd ffipg_2/ffi_1/nand_1/b 0.57fF
C607 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C608 gnd ffipg_0/ffi_1/inv_1/op 1.85fF
C609 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C610 sumffo_2/xor_0/inv_1/op gnd 0.35fF
C611 nor_0/w_0_0# gnd 0.46fF
C612 ffipg_7/ffi_0/q ffipg_7/ffi_0/qbar 0.32fF
C613 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/b 0.32fF
C614 ffipg_6/ffi_1/nand_3/w_0_0# ffipg_6/ffi_1/nand_3/a 0.06fF
C615 gnd ffipg_5/pggen_0/nand_0/w_0_0# 0.10fF
C616 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C617 ffipg_4/ffi_0/nand_3/w_0_0# ffipg_4/ffi_0/nand_3/a 0.06fF
C618 ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C619 gnd ffipg_1/ffi_1/nand_3/a 0.33fF
C620 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/nand_1/b 0.06fF
C621 inv_3/in nor_2/b 0.04fF
C622 cla_2/l cla_2/p0 0.16fF
C623 ffipg_6/ffi_1/q ffipg_6/ffi_1/qbar 0.32fF
C624 gnd sumffo_3/ffo_0/nand_1/w_0_0# 0.10fF
C625 ffipg_6/ffi_1/nand_1/a ffipg_6/ffi_1/nand_1/b 0.31fF
C626 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C627 sumffo_2/xor_0/w_n3_4# ffipg_2/k 0.06fF
C628 gnd ffipg_2/ffi_1/nand_1/a 0.44fF
C629 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a 0.13fF
C630 cla_0/n inv_5/in 0.13fF
C631 cla_0/g0 nand_2/b 0.13fF
C632 ffipg_6/pggen_0/xor_0/w_n3_4# ffipg_6/k 0.02fF
C633 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_1/b 0.31fF
C634 ffi_1/nand_1/a ffi_1/nand_1/b 0.31fF
C635 gnd ffo_0/nand_1/b 0.57fF
C636 ffipg_4/ffi_0/nand_1/a ffipg_4/ffi_0/nand_0/w_0_0# 0.04fF
C637 ffipg_1/ffi_0/inv_0/op y2in 0.04fF
C638 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/inv_1/w_0_6# 0.04fF
C639 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C640 ffi_0/q sumffo_3/ffo_0/d 0.16fF
C641 ffipg_5/ffi_0/nand_5/w_0_0# ffipg_5/ffi_0/nand_7/a 0.04fF
C642 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/nand_7/a 0.04fF
C643 ffi_1/nand_5/w_0_0# ffi_1/nand_7/a 0.04fF
C644 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a 0.31fF
C645 cla_1/p0 ffipg_1/ffi_1/q 0.22fF
C646 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C647 nor_3/w_0_0# nor_3/b 0.06fF
C648 sumffo_3/ffo_0/nand_7/a z4o 0.00fF
C649 sumffo_2/xor_0/w_n3_4# sumffo_2/ffo_0/d 0.02fF
C650 sumffo_0/ffo_0/nand_1/b gnd 0.57fF
C651 ffipg_7/ffi_1/inv_1/op ffipg_7/ffi_1/nand_1/b 0.45fF
C652 ffipg_6/ffi_1/inv_1/op ffipg_6/ffi_1/inv_1/w_0_6# 0.04fF
C653 ffipg_6/ffi_0/nand_3/a gnd 0.33fF
C654 gnd ffipg_4/ffi_1/nand_3/b 0.74fF
C655 gnd ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C656 gnd nor_3/w_0_0# 0.15fF
C657 gnd sumffo_1/ffo_0/nand_1/a 0.44fF
C658 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C659 ffi_0/q sumffo_3/xor_0/a_10_10# 0.04fF
C660 clk ffi_0/inv_1/w_0_6# 0.06fF
C661 gnd nor_0/b 0.74fF
C662 gnd ffipg_2/ffi_1/nand_3/b 0.74fF
C663 ffipg_0/ffi_1/q ffipg_0/ffi_0/q 0.73fF
C664 sumffo_2/ffo_0/nand_7/a z3o 0.00fF
C665 cla_2/g1 gnd 0.65fF
C666 ffipg_4/pggen_0/xor_0/w_n3_4# ffipg_4/pggen_0/xor_0/a_10_10# 0.16fF
C667 ffipg_4/ffi_1/q ffipg_4/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C668 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_1/b 0.45fF
C669 gnd ffo_0/nand_4/w_0_0# 0.10fF
C670 cla_0/l cla_0/n 0.19fF
C671 ffipg_7/ffi_1/inv_1/op x4in 0.01fF
C672 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# 0.04fF
C673 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a 0.13fF
C674 ffipg_1/ffi_0/nand_0/w_0_0# ffipg_1/ffi_0/nand_1/a 0.04fF
C675 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C676 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C677 ffi_1/nand_4/w_0_0# ffi_1/nand_3/b 0.06fF
C678 ffo_0/d inv_9/in 0.04fF
C679 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C680 sumffo_0/ffo_0/nand_4/w_0_0# gnd 0.10fF
C681 ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_1/inv_1/op 0.75fF
C682 ffipg_7/ffi_1/nand_0/w_0_0# clk 0.06fF
C683 ffipg_4/ffi_0/nand_5/w_0_0# ffipg_4/ffi_0/nand_7/a 0.04fF
C684 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_7/a 0.04fF
C685 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C686 ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_7/w_0_0# 0.04fF
C687 gnd ffi_0/nand_4/w_0_0# 0.10fF
C688 ffipg_0/ffi_0/nand_7/w_0_0# ffipg_0/ffi_0/nand_7/a 0.06fF
C689 inv_8/w_0_6# nor_4/a 0.03fF
C690 nor_2/w_0_0# inv_4/in 0.11fF
C691 gnd sumffo_1/xor_0/a_10_10# 0.93fF
C692 ffipg_7/ffi_1/inv_0/op gnd 0.27fF
C693 gnd ffipg_5/ffi_1/inv_0/op 0.27fF
C694 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C695 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/nand_7/a 0.04fF
C696 clk ffipg_2/ffi_0/nand_3/a 0.13fF
C697 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C698 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C699 ffipg_6/ffi_0/q ffipg_6/ffi_0/qbar 0.32fF
C700 ffipg_3/ffi_0/inv_0/op ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C701 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/inv_1/op 0.13fF
C702 ffipg_4/ffi_0/nand_3/b ffipg_4/ffi_0/nand_1/b 0.32fF
C703 sumffo_2/xor_0/w_n3_4# ffi_0/q 0.00fF
C704 ffipg_4/ffi_1/q ffipg_4/k 0.46fF
C705 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C706 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/nand_6/a 0.04fF
C707 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C708 ffipg_6/ffi_0/nand_3/w_0_0# ffipg_6/ffi_0/nand_3/a 0.06fF
C709 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C710 clk ffipg_4/ffi_1/nand_3/a 0.13fF
C711 gnd ffipg_4/ffi_0/inv_0/w_0_6# 0.06fF
C712 ffipg_5/ffi_0/q ffipg_5/ffi_0/qbar 0.32fF
C713 ffipg_5/ffi_0/nand_3/a ffipg_5/ffi_0/nand_3/b 0.31fF
C714 gnd ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C715 gnd ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C716 ffipg_1/ffi_1/nand_6/w_0_0# ffipg_1/ffi_1/qbar 0.04fF
C717 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C718 gnd ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C719 cla_2/l inv_7/w_0_6# 0.06fF
C720 gnd ffipg_3/ffi_0/nand_0/a_13_n26# 0.01fF
C721 gnd ffipg_1/ffi_1/nand_6/a 0.37fF
C722 gnd y2in 0.44fF
C723 ffipg_0/ffi_0/nand_1/w_0_0# ffipg_0/ffi_0/nand_1/a 0.06fF
C724 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C725 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/sbar 0.04fF
C726 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_1/w_0_6# 0.03fF
C727 ffipg_7/ffi_0/nand_5/w_0_0# ffipg_7/ffi_0/inv_1/op 0.06fF
C728 gnd ffipg_4/ffi_0/nand_0/w_0_0# 0.10fF
C729 gnd ffipg_5/ffi_0/nand_2/w_0_0# 0.10fF
C730 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar 0.32fF
C731 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C732 clk sumffo_3/ffo_0/nand_6/a 0.13fF
C733 ffipg_6/ffi_0/q ffipg_6/pggen_0/nor_0/w_0_0# 0.06fF
C734 ffipg_6/ffi_1/q ffipg_6/pggen_0/xor_0/inv_0/op 0.27fF
C735 ffi_0/nand_6/w_0_0# ffi_0/nand_6/a 0.06fF
C736 ffi_0/q inv_0/in 0.07fF
C737 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C738 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/ffi_0/q 0.06fF
C739 sumffo_3/xor_0/inv_0/op inv_4/op 0.27fF
C740 ffipg_7/ffi_0/nand_3/a gnd 0.33fF
C741 ffipg_6/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C742 ffipg_5/g ffipg_5/pggen_0/nand_0/w_0_0# 0.04fF
C743 gnd ffipg_4/ffi_0/inv_1/op 1.85fF
C744 gnd ffipg_5/ffi_1/nand_1/a 0.44fF
C745 ffipg_3/k ffipg_3/ffi_0/q 0.07fF
C746 ffi_1/nand_7/w_0_0# ffi_1/nand_7/a 0.06fF
C747 ffi_1/qbar cinq 0.32fF
C748 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a 0.13fF
C749 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/nand_7/a 0.06fF
C750 gnd ffipg_0/ffi_0/inv_1/op 1.85fF
C751 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_0/b 0.40fF
C752 ffipg_7/ffi_1/qbar ffipg_7/ffi_1/nand_7/a 0.31fF
C753 ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/inv_1/op 0.33fF
C754 ffi_0/nand_3/a ffi_0/nand_3/b 0.31fF
C755 ffipg_0/k ffi_0/q 0.19fF
C756 ffipg_7/ffi_0/nand_0/w_0_0# clk 0.06fF
C757 ffi_0/q sumffo_1/xor_0/inv_0/op 0.06fF
C758 ffipg_4/ffi_1/nand_1/a ffipg_4/ffi_1/nand_1/b 0.31fF
C759 clk ffipg_4/ffi_0/inv_1/w_0_6# 0.06fF
C760 clk ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C761 sumffo_1/ffo_0/nand_6/w_0_0# z2o 0.06fF
C762 cla_1/p0 nor_0/a 0.24fF
C763 gnd ffipg_3/ffi_0/nand_0/w_0_0# 0.10fF
C764 gnd ffipg_2/ffi_1/nand_6/w_0_0# 0.10fF
C765 gnd ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C766 ffo_0/nand_1/a ffo_0/nand_0/w_0_0# 0.04fF
C767 sumffo_0/ffo_0/nand_2/w_0_0# gnd 0.10fF
C768 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/nand_7/a 0.06fF
C769 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/b 0.31fF
C770 clk ffi_0/nand_3/a 0.13fF
C771 ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C772 ffipg_6/pggen_0/nand_0/w_0_0# ffipg_6/ffi_1/q 0.06fF
C773 ffipg_4/ffi_0/nand_6/a ffipg_4/ffi_0/qbar 0.00fF
C774 ffipg_4/ffi_0/q ffipg_4/pggen_0/nor_0/w_0_0# 0.06fF
C775 ffipg_5/ffi_1/nand_1/w_0_0# ffipg_5/ffi_1/nand_1/b 0.06fF
C776 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/a 0.06fF
C777 ffi_0/inv_0/op cinin 0.04fF
C778 gnd ffipg_4/ffi_1/inv_0/w_0_6# 0.06fF
C779 gnd ffipg_2/ffi_0/inv_0/op 0.27fF
C780 ffipg_7/ffi_0/nand_3/b gnd 0.74fF
C781 ffipg_6/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C782 ffipg_6/ffi_0/nand_5/w_0_0# ffipg_6/ffi_0/inv_1/op 0.06fF
C783 gnd ffipg_1/ffi_1/nand_0/a_13_n26# 0.01fF
C784 gnd ffi_0/nand_1/b 0.57fF
C785 ffi_0/nand_1/a ffi_0/nand_1/b 0.31fF
C786 ffi_1/nand_6/a ffi_1/qbar 0.00fF
C787 ffi_0/q sumffo_0/xor_0/a_10_10# 0.12fF
C788 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_3/b 0.04fF
C789 ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_7/w_0_0# 0.04fF
C790 inv_4/op nor_2/w_0_0# 0.03fF
C791 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/ffo_0/nand_6/a 0.06fF
C792 gnd sumffo_1/ffo_0/d 0.41fF
C793 ffipg_7/ffi_0/nand_7/w_0_0# gnd 0.10fF
C794 ffipg_7/ffi_0/inv_0/op clk 0.32fF
C795 ffipg_7/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C796 ffipg_6/ffi_0/nand_5/w_0_0# ffipg_6/ffi_0/nand_7/a 0.04fF
C797 gnd ffipg_3/ffi_1/nand_1/a 0.44fF
C798 gnd inv_9/in 0.33fF
C799 gnd ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C800 gnd ffipg_3/ffi_0/q 3.00fF
C801 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar 0.32fF
C802 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/b 0.31fF
C803 gnd ffipg_0/ffi_1/qbar 0.67fF
C804 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C805 gnd sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C806 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C807 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/nand_1/a 0.04fF
C808 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/inv_0/w_0_6# 0.03fF
C809 sumffo_0/ffo_0/nand_1/w_0_0# gnd 0.10fF
C810 ffipg_7/ffi_0/nand_3/w_0_0# ffipg_7/ffi_0/nand_1/b 0.04fF
C811 ffipg_5/ffi_1/nand_5/w_0_0# ffipg_5/ffi_1/nand_7/a 0.04fF
C812 ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/nand_1/b 0.32fF
C813 ffipg_5/ffi_0/nand_4/w_0_0# ffipg_5/ffi_0/nand_6/a 0.04fF
C814 ffipg_5/ffi_1/q ffipg_5/p 0.22fF
C815 ffi_1/nand_1/b ffi_1/nand_3/b 0.32fF
C816 gnd ffipg_4/ffi_1/nand_2/w_0_0# 0.10fF
C817 ffipg_5/ffi_1/q ffipg_5/pggen_0/xor_0/w_n3_4# 0.06fF
C818 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C819 ffipg_7/ffi_1/nand_3/w_0_0# ffipg_7/ffi_1/nand_1/b 0.04fF
C820 ffipg_7/ffi_0/nand_1/a clk 0.13fF
C821 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C822 gnd ffipg_4/ffi_1/inv_0/op 0.27fF
C823 gnd ffipg_4/pggen_0/xor_0/inv_0/op 0.32fF
C824 ffipg_4/ffi_0/q ffipg_4/g 0.13fF
C825 ffipg_3/ffi_1/nand_7/w_0_0# ffipg_3/ffi_1/nand_7/a 0.06fF
C826 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/ffi_0/q 0.23fF
C827 clk ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C828 gnd ffipg_1/ffi_0/nand_6/a 0.37fF
C829 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_3/b 0.04fF
C830 ffipg_0/ffi_1/nand_2/w_0_0# ffipg_0/ffi_1/nand_3/a 0.04fF
C831 inv_2/w_0_6# nor_1/b 0.03fF
C832 gnd sumffo_2/ffo_0/nand_4/w_0_0# 0.10fF
C833 cla_1/inv_0/op gnd 0.27fF
C834 cla_0/l ffipg_2/k 0.10fF
C835 ffipg_7/ffi_0/nand_0/w_0_0# ffipg_7/ffi_0/inv_0/op 0.06fF
C836 ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_7/a 0.00fF
C837 gnd ffipg_3/ffi_0/nand_2/w_0_0# 0.10fF
C838 clk ffipg_2/ffi_0/inv_1/op 0.07fF
C839 gnd ffo_0/qbar 0.62fF
C840 gnd ffipg_3/ffi_1/qbar 0.67fF
C841 ffipg_1/pggen_0/nand_0/w_0_0# ffipg_1/ffi_1/q 0.06fF
C842 gnd ffipg_0/ffi_1/nand_1/b 0.57fF
C843 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C844 ffipg_6/ffi_0/nand_1/w_0_0# ffipg_6/ffi_0/nand_1/a 0.06fF
C845 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/w_0_0# 0.04fF
C846 ffipg_4/ffi_1/nand_1/w_0_0# ffipg_4/ffi_1/nand_1/a 0.06fF
C847 ffipg_5/ffi_1/q ffipg_5/ffi_0/q 0.73fF
C848 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/qbar 0.00fF
C849 ffi_0/q sumffo_3/xor_0/a_38_n43# 0.01fF
C850 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b 0.32fF
C851 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a 0.00fF
C852 ffipg_7/ffi_0/nand_0/w_0_0# ffipg_7/ffi_0/nand_1/a 0.04fF
C853 ffipg_5/ffi_0/qbar ffipg_5/ffi_0/nand_7/w_0_0# 0.06fF
C854 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/qbar 0.00fF
C855 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C856 ffi_0/nand_1/w_0_0# ffi_0/nand_3/b 0.04fF
C857 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C858 ffipg_1/ffi_1/inv_0/op x2in 0.04fF
C859 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_1/b 0.45fF
C860 ffipg_0/ffi_1/inv_0/op ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C861 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/inv_1/op 0.06fF
C862 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/a 0.06fF
C863 sumffo_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C864 inv_5/w_0_6# inv_5/in 0.10fF
C865 ffipg_7/ffi_1/inv_0/op ffipg_7/ffi_1/inv_0/w_0_6# 0.03fF
C866 ffipg_7/ffi_1/inv_1/op ffipg_7/ffi_1/nand_6/a 0.13fF
C867 ffipg_6/ffi_0/nand_4/w_0_0# gnd 0.10fF
C868 clk sumffo_2/ffo_0/nand_1/b 0.45fF
C869 clk ffipg_3/ffi_0/nand_3/a 0.13fF
C870 gnd ffi_1/nand_3/w_0_0# 0.11fF
C871 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/b 0.31fF
C872 nor_2/b inv_3/w_0_6# 0.03fF
C873 gnd sumffo_3/ffo_0/nand_7/a 0.33fF
C874 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C875 ffipg_6/pggen_0/nor_0/a_13_6# ffipg_6/k 0.01fF
C876 ffipg_5/ffi_0/nand_1/w_0_0# ffipg_5/ffi_0/nand_3/b 0.04fF
C877 ffipg_2/ffi_1/nand_2/w_0_0# x3in 0.06fF
C878 ffi_1/nand_1/a ffi_1/nand_1/w_0_0# 0.06fF
C879 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C880 gnd ffipg_2/ffi_0/nand_3/w_0_0# 0.11fF
C881 ffipg_6/ffi_0/nand_1/a ffipg_6/ffi_0/nand_1/b 0.31fF
C882 ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_6/w_0_0# 0.06fF
C883 ffipg_1/ffi_1/nand_6/w_0_0# ffipg_1/ffi_1/nand_6/a 0.06fF
C884 ffipg_5/pggen_0/nor_0/w_0_0# ffipg_5/k 0.21fF
C885 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/pggen_0/xor_0/inv_1/op 0.08fF
C886 cla_2/p0 ffipg_2/k 0.05fF
C887 ffipg_6/ffi_1/qbar ffipg_6/ffi_1/nand_6/w_0_0# 0.04fF
C888 gnd ffipg_4/ffi_0/nand_2/w_0_0# 0.10fF
C889 ffipg_5/ffi_1/qbar ffipg_5/ffi_1/nand_7/w_0_0# 0.06fF
C890 gnd ffipg_5/ffi_0/nand_5/w_0_0# 0.10fF
C891 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C892 gnd ffi_1/inv_1/op 1.89fF
C893 gnd ffipg_1/ffi_1/q 2.24fF
C894 gnd ffipg_0/ffi_0/nand_2/w_0_0# 0.10fF
C895 inv_6/in nor_3/b 0.16fF
C896 cla_0/l cla_0/inv_0/op 0.35fF
C897 ffipg_6/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C898 gnd sumffo_3/ffo_0/nand_4/w_0_0# 0.10fF
C899 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_1/w_0_6# 0.03fF
C900 cla_2/nor_0/w_0_0# gnd 0.31fF
C901 gnd ffipg_3/ffi_1/nand_3/a 0.33fF
C902 gnd inv_6/in 0.33fF
C903 ffipg_4/ffi_0/nand_1/a ffipg_4/ffi_0/nand_1/b 0.31fF
C904 gnd ffipg_3/ffi_1/nand_3/w_0_0# 0.11fF
C905 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C906 clk ffipg_0/ffi_1/inv_1/op 0.07fF
C907 nor_2/w_0_0# cla_1/n 0.06fF
C908 sumffo_0/xor_0/inv_0/w_0_6# ffipg_0/k 0.06fF
C909 inv_2/in inv_2/w_0_6# 0.10fF
C910 ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/nand_1/b 0.31fF
C911 ffipg_6/pggen_0/nor_0/w_0_0# ffipg_6/p 0.05fF
C912 ffipg_6/pggen_0/xor_0/inv_1/op ffipg_6/pggen_0/xor_0/w_n3_4# 0.06fF
C913 ffi_0/nand_1/b ffi_0/nand_3/w_0_0# 0.04fF
C914 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a 0.00fF
C915 gnd ffo_0/nand_3/b 0.74fF
C916 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/ffi_1/q 0.27fF
C917 ffipg_6/ffi_1/inv_0/op ffipg_6/ffi_1/nand_0/w_0_0# 0.06fF
C918 ffipg_6/ffi_0/nand_6/w_0_0# ffipg_6/ffi_0/qbar 0.04fF
C919 ffipg_4/ffi_0/nand_5/w_0_0# ffipg_4/ffi_0/inv_1/op 0.06fF
C920 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C921 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C922 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op 0.06fF
C923 ffipg_6/ffi_1/inv_1/op ffipg_6/ffi_1/nand_3/b 0.33fF
C924 ffipg_6/ffi_1/nand_1/a ffipg_6/ffi_1/nand_0/w_0_0# 0.04fF
C925 gnd ffipg_1/ffi_0/nand_0/a_13_n26# 0.01fF
C926 clk ffipg_1/ffi_1/nand_3/a 0.13fF
C927 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a 0.00fF
C928 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C929 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C930 sumffo_0/ffo_0/nand_3/b gnd 0.74fF
C931 cla_2/p1 cla_2/inv_0/in 0.02fF
C932 cla_0/l ffi_0/q 0.33fF
C933 gnd sumffo_1/ffo_0/nand_2/a_13_n26# 0.01fF
C934 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C935 sumffo_1/sbar sumffo_1/ffo_0/nand_7/a 0.31fF
C936 ffipg_6/ffi_1/inv_1/op gnd 1.85fF
C937 gnd ffipg_5/ffi_0/nand_1/a 0.44fF
C938 ffipg_5/ffi_1/nand_4/w_0_0# ffipg_5/ffi_1/nand_3/b 0.06fF
C939 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C940 clk ffipg_2/ffi_1/nand_1/a 0.13fF
C941 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C942 inv_8/in nor_4/a 0.04fF
C943 sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# 0.02fF
C944 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/inv_0/w_0_6# 0.03fF
C945 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C946 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/w_0_0# 0.04fF
C947 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/inv_1/op 0.06fF
C948 x4in ffipg_3/ffi_1/inv_1/op 0.01fF
C949 ffipg_3/ffi_1/nand_2/w_0_0# x4in 0.06fF
C950 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C951 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/a 0.06fF
C952 gnd ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C953 inv_7/op inv_7/w_0_6# 0.03fF
C954 clk ffo_0/nand_1/b 0.45fF
C955 gnd inv_2/w_0_6# 0.17fF
C956 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/inv_1/op 0.33fF
C957 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/w_0_0# 0.06fF
C958 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C959 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_1/q 0.06fF
C960 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C961 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C962 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C963 clk sumffo_0/ffo_0/nand_1/b 0.45fF
C964 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C965 cla_0/nand_0/w_0_0# cla_0/l 0.06fF
C966 ffipg_6/ffi_0/nand_3/a clk 0.13fF
C967 cla_0/g0 ffi_0/q 0.08fF
C968 ffipg_7/ffi_0/inv_1/w_0_6# gnd 0.06fF
C969 ffipg_7/ffi_1/q ffipg_7/pggen_0/xor_0/inv_1/op 0.06fF
C970 ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_0/inv_1/w_0_6# 0.04fF
C971 ffipg_5/ffi_0/inv_0/op ffipg_5/ffi_0/inv_0/w_0_6# 0.03fF
C972 clk ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C973 gnd ffipg_3/ffi_0/nand_6/a 0.37fF
C974 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C975 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar 0.32fF
C976 ffipg_0/ffi_1/nand_2/w_0_0# x1in 0.06fF
C977 ffipg_1/ffi_1/nand_3/w_0_0# ffipg_1/ffi_1/nand_1/b 0.04fF
C978 ffipg_6/ffi_0/nand_1/a ffipg_6/ffi_0/nand_0/w_0_0# 0.04fF
C979 x1in ffipg_4/ffi_1/inv_1/op 0.01fF
C980 ffipg_4/ffi_1/nand_3/a ffipg_4/ffi_1/nand_3/b 0.31fF
C981 ffipg_4/pggen_0/xor_0/inv_0/op ffipg_4/pggen_0/xor_0/inv_1/op 0.08fF
C982 cla_0/l cla_1/l 0.08fF
C983 ffipg_7/ffi_1/inv_1/op ffipg_7/ffi_1/inv_1/w_0_6# 0.04fF
C984 ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/inv_0/op 0.20fF
C985 ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/nand_1/b 0.13fF
C986 ffipg_4/ffi_0/qbar ffipg_4/ffi_0/nand_7/w_0_0# 0.06fF
C987 ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_7/w_0_0# 0.04fF
C988 clk ffo_0/nand_4/w_0_0# 0.06fF
C989 ffipg_7/ffi_1/nand_0/w_0_0# ffipg_7/ffi_1/inv_0/op 0.06fF
C990 ffipg_7/ffi_0/nand_3/w_0_0# gnd 0.11fF
C991 gnd ffipg_4/ffi_0/nand_1/b 0.57fF
C992 gnd ffipg_4/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C993 x2in ffipg_5/ffi_1/nand_2/w_0_0# 0.06fF
C994 gnd ffi_1/inv_1/w_0_6# 0.06fF
C995 gnd ffipg_0/ffi_0/nand_1/b 0.57fF
C996 cla_0/n nor_1/b 0.36fF
C997 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C998 ffipg_7/ffi_1/q gnd 2.24fF
C999 nand_2/b inv_2/in 0.34fF
C1000 ffipg_5/ffi_0/nand_3/b ffipg_5/ffi_0/nand_1/b 0.32fF
C1001 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_1/q 0.06fF
C1002 ffi_0/nand_4/w_0_0# ffi_0/nand_3/b 0.06fF
C1003 ffi_1/nand_5/w_0_0# ffi_1/inv_1/op 0.06fF
C1004 sumffo_0/ffo_0/nand_4/w_0_0# clk 0.06fF
C1005 cla_2/l nor_3/b 0.10fF
C1006 gnd ffipg_0/ffi_1/nand_3/w_0_0# 0.11fF
C1007 ffo_0/nand_1/a ffo_0/nand_1/w_0_0# 0.06fF
C1008 gnd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C1009 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C1010 gnd nor_0/a 0.53fF
C1011 gnd ffipg_4/ffi_1/nand_1/b 0.57fF
C1012 gnd ffipg_2/ffi_0/nand_1/b 0.57fF
C1013 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C1014 cla_0/g0 ffipg_1/k 0.06fF
C1015 gnd ffipg_2/ffi_1/nand_6/a 0.37fF
C1016 gnd ffipg_1/ffi_0/nand_3/a 0.33fF
C1017 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_1/b 0.31fF
C1018 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_0/op 0.08fF
C1019 cla_2/l gnd 0.57fF
C1020 ffipg_4/ffi_0/nand_1/w_0_0# ffipg_4/ffi_0/nand_3/b 0.04fF
C1021 clk ffipg_5/ffi_1/inv_0/op 0.32fF
C1022 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/qbar 0.00fF
C1023 ffipg_7/ffi_1/inv_0/op clk 0.32fF
C1024 ffipg_6/pggen_0/nand_0/w_0_0# ffipg_6/ffi_0/q 0.06fF
C1025 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_1/w_0_6# 0.03fF
C1026 ffipg_7/pggen_0/nor_0/w_0_0# gnd 0.11fF
C1027 ffipg_6/ffi_0/nand_1/w_0_0# ffipg_6/ffi_0/nand_3/b 0.04fF
C1028 ffipg_6/ffi_0/nand_4/w_0_0# ffipg_6/ffi_0/nand_6/a 0.04fF
C1029 gnd ffipg_5/ffi_1/nand_5/w_0_0# 0.10fF
C1030 gnd ffi_1/inv_0/op 0.27fF
C1031 gnd ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C1032 gnd sumffo_2/ffo_0/nand_1/a 0.33fF
C1033 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C1034 cla_1/l cla_2/p0 0.02fF
C1035 cla_1/p0 ffipg_2/k 0.06fF
C1036 gnd ffo_0/inv_0/w_0_6# 0.07fF
C1037 gnd nand_2/b 1.93fF
C1038 gnd ffipg_4/ffi_0/qbar 0.67fF
C1039 gnd ffipg_5/pggen_0/nor_0/w_0_0# 0.11fF
C1040 clk ffipg_4/ffi_0/nand_0/w_0_0# 0.06fF
C1041 clk ffipg_5/ffi_0/nand_2/w_0_0# 0.06fF
C1042 ffipg_2/ffi_1/nand_2/w_0_0# ffipg_2/ffi_1/nand_3/a 0.04fF
C1043 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.32fF
C1044 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C1045 clk y2in 1.36fF
C1046 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.32fF
C1047 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/inv_1/op 0.33fF
C1048 sumffo_0/xor_0/inv_0/op ffi_0/q 0.20fF
C1049 ffipg_6/ffi_0/inv_0/op ffipg_6/ffi_0/nand_0/w_0_0# 0.06fF
C1050 y1in ffipg_4/ffi_0/inv_0/op 0.04fF
C1051 ffi_1/nand_1/w_0_0# ffi_1/nand_3/b 0.04fF
C1052 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/w_0_0# 0.06fF
C1053 ffo_0/qbar couto 0.32fF
C1054 x3in ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C1055 ffipg_3/ffi_1/inv_0/op ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1056 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C1057 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/nand_1/b 0.06fF
C1058 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.35fF
C1059 ffipg_0/ffi_1/nand_4/w_0_0# ffipg_0/ffi_1/inv_1/op 0.06fF
C1060 gnd nor_4/b 0.25fF
C1061 ffipg_7/ffi_0/nand_3/a clk 0.13fF
C1062 ffipg_6/ffi_1/inv_0/w_0_6# gnd 0.06fF
C1063 ffipg_6/ffi_0/inv_0/w_0_6# y3in 0.06fF
C1064 ffipg_7/ffi_1/nand_6/w_0_0# ffipg_7/ffi_1/nand_6/a 0.06fF
C1065 ffipg_6/ffi_0/nand_3/b ffipg_6/ffi_0/nand_1/b 0.32fF
C1066 clk ffipg_4/ffi_0/inv_1/op 0.07fF
C1067 ffipg_4/ffi_0/nand_3/w_0_0# ffipg_4/ffi_0/nand_3/b 0.06fF
C1068 clk ffipg_5/ffi_1/nand_1/a 0.13fF
C1069 gnd ffi_1/nand_6/w_0_0# 0.10fF
C1070 ffipg_2/ffi_1/nand_4/w_0_0# ffipg_2/ffi_1/nand_6/a 0.04fF
C1071 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_1/b 0.31fF
C1072 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1073 clk ffipg_0/ffi_0/inv_1/op 0.07fF
C1074 ffipg_3/k cla_0/n 0.06fF
C1075 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C1076 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C1077 ffipg_4/ffi_1/q ffipg_4/ffi_1/nand_7/a 0.00fF
C1078 gnd y4in 0.44fF
C1079 gnd ffipg_4/ffi_1/nand_1/w_0_0# 0.10fF
C1080 clk ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C1081 gnd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C1082 gnd sumffo_3/ffo_0/inv_0/w_0_6# 0.07fF
C1083 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C1084 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C1085 ffipg_6/ffi_0/inv_1/op y3in 0.01fF
C1086 ffi_0/nand_1/b ffi_0/nand_3/b 0.32fF
C1087 ffi_1/inv_0/w_0_6# cinin 0.06fF
C1088 clk ffipg_2/ffi_0/inv_0/op 0.32fF
C1089 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/k 0.06fF
C1090 ffipg_7/ffi_0/nand_1/b ffipg_7/ffi_0/nand_7/a 0.13fF
C1091 gnd ffipg_4/ffi_1/q 2.24fF
C1092 ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_0/inv_1/w_0_6# 0.04fF
C1093 ffipg_5/ffi_0/qbar ffipg_5/ffi_0/nand_7/a 0.31fF
C1094 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C1095 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C1096 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_7/a 0.04fF
C1097 sumffo_0/ffo_0/nand_7/w_0_0# z1o 0.04fF
C1098 gnd sumffo_1/sbar 0.62fF
C1099 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C1100 ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_0/inv_1/w_0_6# 0.04fF
C1101 gnd ffipg_5/ffi_0/nand_3/a 0.33fF
C1102 gnd ffipg_2/ffi_1/nand_0/w_0_0# 0.10fF
C1103 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/inv_1/w_0_6# 0.04fF
C1104 ffi_0/q sumffo_2/xor_0/a_38_n43# 0.01fF
C1105 clk sumffo_1/ffo_0/d 0.04fF
C1106 clk ffipg_3/ffi_1/nand_1/a 0.13fF
C1107 gnd ffipg_4/pggen_0/nand_0/w_0_0# 0.10fF
C1108 gnd ffipg_5/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1109 gnd ffipg_2/ffi_0/nand_3/b 0.74fF
C1110 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C1111 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C1112 cla_0/l ffipg_1/ffi_0/q 0.13fF
C1113 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1114 sumffo_3/ffo_0/d sumffo_3/xor_0/a_10_10# 0.45fF
C1115 clk sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C1116 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1117 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C1118 cla_2/inv_0/op gnd 0.27fF
C1119 ffipg_7/ffi_1/nand_5/w_0_0# gnd 0.10fF
C1120 ffipg_4/ffi_1/q p1 0.22fF
C1121 gnd cla_0/n 0.87fF
C1122 ffipg_6/ffi_1/inv_0/op gnd 0.27fF
C1123 ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_6/a 0.31fF
C1124 clk ffipg_4/ffi_1/nand_2/w_0_0# 0.06fF
C1125 ffipg_6/ffi_1/nand_1/a ffipg_6/ffi_1/nand_3/b 0.00fF
C1126 ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/nand_6/w_0_0# 0.06fF
C1127 ffipg_6/ffi_1/nand_1/a gnd 0.44fF
C1128 ffipg_4/ffi_1/nand_3/a ffipg_4/ffi_1/nand_2/w_0_0# 0.04fF
C1129 clk ffipg_4/ffi_1/inv_0/op 0.32fF
C1130 ffipg_4/pggen_0/nand_0/w_0_0# p1 0.24fF
C1131 ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/inv_0/op 0.20fF
C1132 ffipg_5/ffi_1/qbar ffipg_5/ffi_1/nand_7/a 0.31fF
C1133 ffipg_5/ffi_0/nand_1/b ffipg_5/ffi_0/nand_7/a 0.13fF
C1134 gnd ffipg_5/ffi_0/inv_1/op 1.85fF
C1135 gnd ffi_1/nand_4/w_0_0# 0.10fF
C1136 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_1/b 0.31fF
C1137 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C1138 gnd z2o 0.80fF
C1139 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1140 clk sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C1141 sumffo_2/ffo_0/nand_3/w_0_0# gnd 0.11fF
C1142 ffipg_4/pggen_0/xor_0/inv_1/w_0_6# ffipg_4/pggen_0/xor_0/inv_1/op 0.03fF
C1143 ffipg_7/k ffipg_7/pggen_0/xor_0/inv_1/op 0.52fF
C1144 ffipg_4/ffi_1/qbar ffipg_4/ffi_1/nand_7/a 0.31fF
C1145 clk ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1146 gnd ffi_0/nand_7/a 0.33fF
C1147 cla_2/p0 ffipg_2/ffi_1/q 0.22fF
C1148 ffipg_6/pggen_0/nor_0/w_0_0# ffipg_6/k 0.21fF
C1149 ffipg_5/ffi_1/nand_5/w_0_0# ffipg_5/ffi_1/inv_1/op 0.06fF
C1150 y3in ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C1151 ffipg_0/ffi_0/nand_1/w_0_0# ffipg_0/ffi_0/nand_3/b 0.04fF
C1152 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# 0.04fF
C1153 ffipg_6/ffi_0/nand_1/a gnd 0.44fF
C1154 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/qbar 0.00fF
C1155 ffipg_4/ffi_0/nand_5/w_0_0# ffipg_4/ffi_0/nand_1/b 0.06fF
C1156 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C1157 cla_0/inv_0/w_0_6# cla_0/inv_0/op 0.03fF
C1158 ffipg_7/k gnd 0.27fF
C1159 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/pggen_0/xor_0/w_n3_4# 0.06fF
C1160 gnd ffipg_4/ffi_1/qbar 0.67fF
C1161 ffipg_5/ffi_1/nand_1/b ffipg_5/ffi_1/nand_7/a 0.13fF
C1162 gnd ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C1163 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b 0.32fF
C1164 ffipg_1/ffi_0/nand_3/w_0_0# ffipg_1/ffi_0/nand_1/b 0.04fF
C1165 nor_0/a ffipg_0/ffi_1/q 0.22fF
C1166 nor_0/w_0_0# nor_0/b 0.06fF
C1167 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/ffo_0/nand_7/a 0.06fF
C1168 sumffo_3/sbar z4o 0.32fF
C1169 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C1170 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C1171 ffi_0/q sumffo_2/xor_0/a_10_10# 0.04fF
C1172 cla_1/p0 ffipg_1/k 0.05fF
C1173 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a 0.00fF
C1174 ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C1175 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C1176 ffipg_7/ffi_1/q ffipg_7/ffi_1/nand_7/a 0.00fF
C1177 ffipg_6/ffi_1/qbar ffipg_6/ffi_1/nand_7/a 0.31fF
C1178 sumffo_3/xor_0/w_n3_4# inv_4/op 0.06fF
C1179 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C1180 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C1181 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C1182 nor_2/b inv_4/in 0.16fF
C1183 nor_1/w_0_0# nor_1/b 0.06fF
C1184 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_0/b 0.40fF
C1185 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C1186 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C1187 cla_0/l cla_2/p1 0.30fF
C1188 cla_1/p0 cla_1/l 0.16fF
C1189 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/a 0.00fF
C1190 gnd x3in 0.44fF
C1191 ffipg_6/pggen_0/nand_0/w_0_0# ffipg_6/p 0.24fF
C1192 ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/a_10_10# 0.12fF
C1193 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/inv_1/op 0.33fF
C1194 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C1195 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_3/b 0.06fF
C1196 inv_7/op inv_7/in 0.04fF
C1197 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C1198 ffipg_7/ffi_1/nand_4/w_0_0# ffipg_7/ffi_1/inv_1/op 0.06fF
C1199 ffipg_4/ffi_0/nand_1/w_0_0# ffipg_4/ffi_0/nand_1/a 0.06fF
C1200 ffi_0/nand_1/b ffi_0/nand_5/w_0_0# 0.06fF
C1201 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C1202 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b 0.32fF
C1203 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a 0.31fF
C1204 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C1205 clk ffipg_4/ffi_0/nand_2/w_0_0# 0.06fF
C1206 ffipg_4/pggen_0/xor_0/w_n3_4# ffipg_4/k 0.02fF
C1207 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_1/b 0.45fF
C1208 clk ffi_1/inv_1/op 0.93fF
C1209 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a 0.00fF
C1210 clk ffipg_0/ffi_0/nand_2/w_0_0# 0.06fF
C1211 gnd ffipg_2/ffi_0/nand_6/a 0.37fF
C1212 clk sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C1213 gnd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C1214 clk ffipg_3/ffi_1/nand_3/a 0.13fF
C1215 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C1216 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C1217 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C1218 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/qbar 0.00fF
C1219 ffi_1/inv_0/op ffi_1/nand_0/w_0_0# 0.06fF
C1220 ffipg_7/ffi_0/nand_5/w_0_0# ffipg_7/ffi_0/nand_1/b 0.06fF
C1221 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/ffo_0/nand_6/a 0.06fF
C1222 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C1223 ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/pggen_0/xor_0/w_n3_4# 0.06fF
C1224 ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_7/a 0.00fF
C1225 ffipg_5/ffi_0/nand_3/a ffipg_5/ffi_0/nand_3/w_0_0# 0.06fF
C1226 ffipg_0/ffi_0/inv_0/op y1in 0.04fF
C1227 clk ffo_0/nand_3/b 0.33fF
C1228 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_6/a 0.04fF
C1229 ffipg_6/ffi_1/nand_2/w_0_0# x3in 0.06fF
C1230 ffipg_6/ffi_0/inv_0/op gnd 0.27fF
C1231 inv_7/op gnd 0.27fF
C1232 ffipg_6/ffi_0/qbar gnd 0.67fF
C1233 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C1234 inv_1/in nor_1/b 0.16fF
C1235 gnd sumffo_3/xor_0/inv_0/op 0.32fF
C1236 cla_2/p0 cla_2/p1 0.24fF
C1237 sumffo_0/ffo_0/nand_3/b clk 0.33fF
C1238 gnd ffipg_0/ffi_1/nand_0/a_13_n26# 0.01fF
C1239 gnd sumffo_2/ffo_0/nand_7/a 0.33fF
C1240 ffipg_7/ffi_0/inv_0/w_0_6# gnd 0.06fF
C1241 ffipg_7/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C1242 ffipg_6/ffi_1/inv_1/op clk 0.07fF
C1243 clk ffipg_5/ffi_0/nand_1/a 0.13fF
C1244 gnd ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C1245 gnd ffipg_5/ffi_0/nand_1/w_0_0# 0.10fF
C1246 ffi_0/nand_1/w_0_0# ffi_0/nand_1/b 0.06fF
C1247 gnd ffi_1/nand_1/b 0.57fF
C1248 gnd ffipg_2/ffi_1/nand_1/w_0_0# 0.10fF
C1249 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C1250 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_1/inv_1/op 0.75fF
C1251 sumffo_0/ffo_0/d gnd 0.41fF
C1252 ffipg_4/ffi_1/q ffipg_4/pggen_0/xor_0/inv_1/op 0.06fF
C1253 ffipg_6/ffi_1/q ffipg_6/ffi_0/q 0.73fF
C1254 ffipg_4/pggen_0/xor_0/a_10_10# ffipg_4/k 0.45fF
C1255 ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_1/inv_1/op 0.75fF
C1256 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C1257 inv_9/in nor_4/w_0_0# 0.11fF
C1258 gnd inv_8/w_0_6# 0.15fF
C1259 ffipg_6/pggen_0/nor_0/w_0_0# gnd 0.11fF
C1260 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C1261 cla_1/nor_0/w_0_0# gnd 0.31fF
C1262 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/ffi_0/q 0.20fF
C1263 ffipg_7/g gnd 0.31fF
C1264 ffipg_6/ffi_0/nand_5/w_0_0# ffipg_6/ffi_0/nand_1/b 0.06fF
C1265 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C1266 gnd cinq 0.80fF
C1267 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C1268 gnd ffipg_0/ffi_1/nand_3/a 0.33fF
C1269 gnd sumffo_3/ffo_0/nand_1/b 0.57fF
C1270 gnd sumffo_1/ffo_0/nand_5/w_0_0# 0.10fF
C1271 ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_7/a 0.00fF
C1272 gnd ffi_1/nand_0/a_13_n26# 0.01fF
C1273 gnd ffipg_0/ffi_0/qbar 0.67fF
C1274 gnd nor_2/w_0_0# 0.15fF
C1275 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_3/b 0.04fF
C1276 gnd ffipg_2/k 0.58fF
C1277 ffipg_7/ffi_0/inv_1/w_0_6# clk 0.06fF
C1278 ffipg_7/ffi_0/nand_7/a gnd 0.37fF
C1279 gnd ffipg_3/ffi_1/nand_3/b 0.74fF
C1280 gnd ffipg_4/ffi_0/nand_1/w_0_0# 0.10fF
C1281 gnd ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C1282 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b 0.32fF
C1283 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_1/a 0.04fF
C1284 sumffo_0/ffo_0/nand_0/w_0_0# gnd 0.10fF
C1285 ffipg_5/ffi_0/q ffipg_5/p 0.03fF
C1286 ffo_0/nand_7/w_0_0# ffo_0/nand_7/a 0.06fF
C1287 ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_6/w_0_0# 0.06fF
C1288 ffipg_3/ffi_0/nand_2/w_0_0# ffipg_3/ffi_0/nand_3/a 0.04fF
C1289 ffipg_5/ffi_1/q ffipg_5/k 0.46fF
C1290 ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/w_n3_4# 0.06fF
C1291 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C1292 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C1293 ffipg_7/k ffipg_7/pggen_0/xor_0/a_10_10# 0.45fF
C1294 gnd sumffo_2/ffo_0/d 0.41fF
C1295 ffipg_7/ffi_1/nand_5/w_0_0# ffipg_7/ffi_1/nand_7/a 0.04fF
C1296 ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1297 gnd ffipg_5/ffi_0/inv_0/w_0_6# 0.06fF
C1298 clk ffi_1/inv_1/w_0_6# 0.06fF
C1299 gnd ffi_1/nand_6/a 0.33fF
C1300 gnd ffipg_1/ffi_1/nand_4/w_0_0# 0.10fF
C1301 ffipg_1/ffi_0/nand_6/w_0_0# ffipg_1/ffi_0/nand_6/a 0.06fF
C1302 gnd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C1303 gnd nor_1/w_0_0# 0.15fF
C1304 ffipg_6/ffi_0/nand_7/w_0_0# gnd 0.10fF
C1305 ffipg_5/ffi_0/inv_0/op ffipg_5/ffi_0/nand_0/w_0_0# 0.06fF
C1306 gnd ffipg_5/ffi_1/inv_0/w_0_6# 0.06fF
C1307 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.32fF
C1308 ffi_1/nand_3/a ffi_1/nand_3/b 0.31fF
C1309 gnd ffipg_2/ffi_1/inv_0/op 0.27fF
C1310 gnd ffipg_1/ffi_0/nand_2/w_0_0# 0.10fF
C1311 clk ffipg_1/ffi_0/nand_3/a 0.13fF
C1312 cla_1/p0 ffipg_1/ffi_0/q 0.03fF
C1313 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C1314 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C1315 ffipg_7/ffi_0/nand_1/w_0_0# ffipg_7/ffi_0/nand_1/b 0.06fF
C1316 ffipg_7/pggen_0/xor_0/inv_1/op ffipg_7/ffi_0/q 0.22fF
C1317 ffi_0/q inv_2/in 0.13fF
C1318 sumffo_0/ffo_0/nand_7/a z1o 0.00fF
C1319 sumffo_0/ffo_0/nand_7/w_0_0# gnd 0.10fF
C1320 cla_0/inv_0/op gnd 0.27fF
C1321 ffipg_7/ffi_0/nand_6/w_0_0# ffipg_7/ffi_0/qbar 0.04fF
C1322 ffipg_6/ffi_0/nand_3/b gnd 0.74fF
C1323 gnd ffipg_4/ffi_0/nand_3/w_0_0# 0.11fF
C1324 ffipg_5/ffi_1/nand_1/w_0_0# ffipg_5/ffi_1/nand_3/b 0.04fF
C1325 gnd ffipg_5/ffi_0/qbar 0.67fF
C1326 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/inv_1/w_0_6# 0.04fF
C1327 clk ffi_1/inv_0/op 0.32fF
C1328 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C1329 gnd ffipg_1/ffi_0/nand_5/w_0_0# 0.10fF
C1330 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_1/b 0.45fF
C1331 inv_5/w_0_6# nor_3/b 0.17fF
C1332 gnd sumffo_1/xor_0/inv_1/op 0.35fF
C1333 gnd inv_5/w_0_6# 0.41fF
C1334 ffipg_7/ffi_0/q gnd 3.00fF
C1335 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b 0.32fF
C1336 ffipg_4/ffi_0/q ffipg_4/ffi_0/qbar 0.32fF
C1337 gnd ffipg_5/ffi_1/qbar 0.67fF
C1338 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C1339 gnd ffi_0/inv_0/w_0_6# 0.06fF
C1340 ffi_1/nand_1/b ffi_1/nand_5/w_0_0# 0.06fF
C1341 gnd ffipg_2/ffi_1/nand_3/a 0.33fF
C1342 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C1343 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C1344 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1345 ffipg_7/ffi_1/inv_1/op gnd 1.85fF
C1346 ffipg_6/ffi_1/nand_5/w_0_0# ffipg_6/ffi_1/inv_1/op 0.06fF
C1347 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/nand_7/a 0.04fF
C1348 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/a 0.31fF
C1349 gnd inv_1/in 0.33fF
C1350 y2in ffipg_5/ffi_0/nand_2/w_0_0# 0.06fF
C1351 ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/nand_4/w_0_0# 0.04fF
C1352 cla_2/p1 ffipg_3/ffi_1/q 0.22fF
C1353 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar 0.32fF
C1354 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C1355 ffi_0/q gnd 2.14fF
C1356 ffipg_7/pggen_0/xor_0/w_n3_4# ffipg_7/pggen_0/xor_0/a_10_10# 0.16fF
C1357 ffipg_5/ffi_0/nand_6/w_0_0# ffipg_5/ffi_0/qbar 0.04fF
C1358 gnd ffipg_5/ffi_0/nand_1/b 0.57fF
C1359 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a 0.13fF
C1360 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C1361 cla_2/g1 ffipg_3/ffi_0/q 0.13fF
C1362 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/inv_1/op 0.33fF
C1363 gnd y1in 0.44fF
C1364 gnd sumffo_3/ffo_0/nand_3/w_0_0# 0.11fF
C1365 ffipg_6/ffi_1/qbar gnd 0.67fF
C1366 ffo_0/nand_6/w_0_0# ffo_0/nand_6/a 0.06fF
C1367 clk y4in 1.28fF
C1368 gnd ffipg_5/ffi_1/nand_1/b 0.57fF
C1369 gnd ffipg_3/ffi_1/nand_5/w_0_0# 0.10fF
C1370 gnd ffi_0/nand_2/w_0_0# 0.10fF
C1371 nor_2/b cla_1/n 0.39fF
C1372 gnd sumffo_3/sbar 0.62fF
C1373 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C1374 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C1375 cla_0/l cla_2/inv_0/in 0.16fF
C1376 ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/k 0.06fF
C1377 ffipg_5/ffi_1/nand_3/w_0_0# ffipg_5/ffi_1/nand_1/b 0.04fF
C1378 ffipg_3/ffi_1/inv_0/op x4in 0.04fF
C1379 gnd inv_3/in 0.47fF
C1380 ffipg_7/ffi_0/nand_5/w_0_0# gnd 0.10fF
C1381 sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# 0.02fF
C1382 ffipg_6/ffi_0/nand_6/a ffipg_6/ffi_0/qbar 0.00fF
C1383 ffipg_1/ffi_0/nand_0/w_0_0# ffipg_1/ffi_0/inv_0/op 0.06fF
C1384 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C1385 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C1386 cla_0/nand_0/w_0_0# gnd 0.10fF
C1387 ffipg_6/ffi_0/nand_3/w_0_0# ffipg_6/ffi_0/nand_3/b 0.06fF
C1388 ffipg_4/ffi_0/q ffipg_4/ffi_1/q 0.73fF
C1389 ffipg_5/ffi_1/nand_6/w_0_0# ffipg_5/ffi_1/qbar 0.04fF
C1390 ffipg_5/ffi_0/inv_1/op ffipg_5/ffi_0/nand_6/a 0.13fF
C1391 gnd ffi_0/nand_0/w_0_0# 0.10fF
C1392 ffi_0/nand_0/w_0_0# ffi_0/nand_1/a 0.04fF
C1393 gnd ffipg_1/ffi_1/nand_2/w_0_0# 0.10fF
C1394 nor_0/a ffipg_0/ffi_0/q 0.03fF
C1395 clk ffipg_5/ffi_0/nand_3/a 0.13fF
C1396 clk ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C1397 gnd ffipg_2/ffi_0/nand_7/w_0_0# 0.10fF
C1398 gnd x1in 0.44fF
C1399 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a 0.13fF
C1400 gnd ffipg_1/k 0.70fF
C1401 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C1402 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C1403 ffipg_4/ffi_0/nand_1/b ffipg_4/ffi_0/nand_7/a 0.13fF
C1404 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a 0.31fF
C1405 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1406 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b 0.32fF
C1407 gnd ffi_0/inv_1/op 1.89fF
C1408 gnd ffipg_2/ffi_1/inv_1/op 1.85fF
C1409 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_1/b 0.45fF
C1410 ffo_0/inv_0/op ffo_0/d 0.04fF
C1411 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C1412 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C1413 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C1414 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C1415 cla_1/l gnd 0.40fF
C1416 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_3/a 0.31fF
C1417 ffipg_6/ffi_1/q ffipg_6/p 0.22fF
C1418 ffipg_4/pggen_0/nor_0/a_13_6# ffipg_4/k 0.01fF
C1419 ffipg_4/ffi_0/q ffipg_4/pggen_0/nand_0/w_0_0# 0.06fF
C1420 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C1421 ffipg_2/k ffipg_2/ffi_0/q 0.07fF
C1422 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.35fF
C1423 gnd ffo_0/nand_3/w_0_0# 0.11fF
C1424 ffipg_7/ffi_0/nand_2/w_0_0# gnd 0.10fF
C1425 ffipg_6/ffi_1/inv_0/op clk 0.32fF
C1426 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# 0.04fF
C1427 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b 0.32fF
C1428 ffipg_6/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C1429 sumffo_0/ffo_0/nand_3/w_0_0# gnd 0.11fF
C1430 ffipg_6/ffi_1/nand_3/w_0_0# ffipg_6/ffi_1/nand_3/b 0.06fF
C1431 ffipg_6/ffi_1/nand_1/a clk 0.13fF
C1432 clk ffipg_5/ffi_0/inv_1/op 0.07fF
C1433 gnd ffipg_5/ffi_1/q 2.24fF
C1434 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C1435 gnd sumffo_2/ffo_0/inv_1/w_0_6# 0.07fF
C1436 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C1437 ffipg_6/ffi_1/nand_3/w_0_0# gnd 0.11fF
C1438 ffipg_4/ffi_1/nand_6/a ffipg_4/ffi_1/inv_1/op 0.13fF
C1439 ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_7/w_0_0# 0.04fF
C1440 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# 0.04fF
C1441 nor_3/w_0_0# inv_6/in 0.11fF
C1442 ffo_0/nand_3/b ffo_0/nand_1/b 0.32fF
C1443 ffipg_7/ffi_1/q ffipg_7/ffi_1/qbar 0.32fF
C1444 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/w_0_0# 0.06fF
C1445 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C1446 ffipg_7/ffi_0/inv_0/op y4in 0.04fF
C1447 ffipg_6/ffi_0/nand_2/w_0_0# y3in 0.06fF
C1448 ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1449 ffipg_4/ffi_0/qbar ffipg_4/ffi_0/nand_7/a 0.31fF
C1450 ffipg_4/ffi_1/q ffipg_4/pggen_0/nor_0/w_0_0# 0.06fF
C1451 ffipg_6/ffi_1/nand_1/w_0_0# ffipg_6/ffi_1/nand_1/a 0.06fF
C1452 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_3/b 0.04fF
C1453 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C1454 ffipg_7/p gnd 0.35fF
C1455 ffipg_6/ffi_0/nand_1/a clk 0.13fF
C1456 gnd sumffo_2/ffo_0/nand_2/w_0_0# 0.10fF
C1457 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d 0.04fF
C1458 ffipg_7/ffi_0/q ffipg_7/pggen_0/xor_0/a_10_10# 0.12fF
C1459 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1460 ffi_1/nand_7/w_0_0# cinq 0.04fF
C1461 sumffo_0/xor_0/inv_1/op ffi_0/q 0.22fF
C1462 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b 0.32fF
C1463 ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/inv_1/op 0.33fF
C1464 ffi_1/nand_2/w_0_0# cinin 0.06fF
C1465 clk ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C1466 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C1467 inv_4/op inv_4/in 0.04fF
C1468 gnd ffipg_3/ffi_0/inv_1/op 1.85fF
C1469 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C1470 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C1471 gnd sumffo_1/ffo_0/nand_3/b 0.74fF
C1472 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/b 0.31fF
C1473 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/b 0.31fF
C1474 ffi_1/nand_1/a ffi_1/nand_3/b 0.00fF
C1475 x2in ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C1476 gnd ffi_1/nand_1/w_0_0# 0.10fF
C1477 gnd ffipg_1/ffi_0/nand_0/w_0_0# 0.10fF
C1478 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C1479 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C1480 sumffo_0/ffo_0/nand_0/b gnd 0.58fF
C1481 ffipg_4/ffi_1/nand_5/w_0_0# ffipg_4/ffi_1/inv_1/op 0.06fF
C1482 ffipg_5/ffi_0/nand_3/w_0_0# ffipg_5/ffi_0/nand_1/b 0.04fF
C1483 clk x3in 1.36fF
C1484 ffipg_6/pggen_0/nand_0/w_0_0# ffipg_6/g 0.04fF
C1485 ffipg_4/ffi_1/inv_0/op ffipg_4/ffi_1/inv_0/w_0_6# 0.03fF
C1486 ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_6/w_0_0# 0.06fF
C1487 x1in ffipg_0/ffi_1/inv_0/op 0.04fF
C1488 nor_0/w_0_0# nor_0/a 0.06fF
C1489 gnd inv_8/in 0.43fF
C1490 ffipg_7/ffi_0/nand_1/w_0_0# gnd 0.10fF
C1491 ffipg_6/pggen_0/xor_0/inv_0/op gnd 0.32fF
C1492 gnd ffo_0/nand_0/w_0_0# 0.10fF
C1493 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/op 0.04fF
C1494 gnd sumffo_2/ffo_0/nand_3/b 0.74fF
C1495 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C1496 cla_2/nand_0/w_0_0# gnd 0.18fF
C1497 ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_0/nand_1/b 0.45fF
C1498 ffipg_4/ffi_1/nand_1/a ffipg_4/ffi_1/nand_0/w_0_0# 0.04fF
C1499 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C1500 x2in ffipg_1/ffi_1/inv_1/op 0.01fF
C1501 ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C1502 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C1503 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C1504 ffipg_5/ffi_1/inv_1/op ffipg_5/ffi_1/nand_1/b 0.45fF
C1505 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C1506 gnd ffipg_3/ffi_1/nand_0/w_0_0# 0.10fF
C1507 nor_4/b nor_4/w_0_0# 0.06fF
C1508 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C1509 ffipg_7/ffi_1/nand_3/w_0_0# gnd 0.11fF
C1510 ffipg_6/ffi_0/nand_1/b ffipg_6/ffi_0/nand_7/a 0.13fF
C1511 gnd ffipg_5/ffi_1/nand_4/w_0_0# 0.10fF
C1512 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/w_0_0# 0.06fF
C1513 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a 0.31fF
C1514 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_1/inv_1/op 0.75fF
C1515 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a 0.31fF
C1516 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_3/b 0.00fF
C1517 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# 0.04fF
C1518 gnd ffipg_0/ffi_1/nand_7/w_0_0# 0.10fF
C1519 sumffo_0/xor_0/w_n3_4# ffi_0/q 0.06fF
C1520 sumffo_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C1521 ffipg_7/ffi_0/nand_4/w_0_0# ffipg_7/ffi_0/inv_1/op 0.06fF
C1522 ffipg_4/g ffipg_4/pggen_0/nand_0/w_0_0# 0.04fF
C1523 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/nand_6/a 0.06fF
C1524 ffipg_4/ffi_0/nand_6/w_0_0# ffipg_4/ffi_0/nand_6/a 0.06fF
C1525 ffipg_6/ffi_0/inv_0/op clk 0.32fF
C1526 ffipg_6/pggen_0/nand_0/w_0_0# gnd 0.10fF
C1527 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1528 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a 0.00fF
C1529 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/inv_1/op 0.33fF
C1530 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C1531 gnd ffo_0/inv_0/op 0.37fF
C1532 nor_0/w_0_0# nand_2/b 0.04fF
C1533 gnd sumffo_1/xor_0/w_n3_4# 0.12fF
C1534 ffipg_6/ffi_0/nand_5/w_0_0# gnd 0.10fF
C1535 ffipg_4/ffi_1/inv_1/op ffipg_4/ffi_1/inv_1/w_0_6# 0.04fF
C1536 ffipg_4/ffi_0/nand_3/a ffipg_4/ffi_0/nand_3/b 0.31fF
C1537 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C1538 gnd ffi_0/nand_7/w_0_0# 0.10fF
C1539 gnd ffipg_2/ffi_1/q 2.24fF
C1540 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/nand_7/a 0.04fF
C1541 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C1542 gnd sumffo_2/ffo_0/nand_3/a 0.33fF
C1543 sumffo_0/ffo_0/d clk 0.25fF
C1544 ffipg_5/ffi_0/nand_4/w_0_0# ffipg_5/ffi_0/inv_1/op 0.06fF
C1545 gnd ffipg_3/ffi_1/nand_7/w_0_0# 0.10fF
C1546 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C1547 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C1548 ffi_0/nand_5/w_0_0# ffi_0/nand_7/a 0.04fF
C1549 gnd x2in 0.44fF
C1550 gnd ffipg_1/ffi_0/q 3.00fF
C1551 sumffo_1/ffo_0/nand_6/a gnd 0.33fF
C1552 ffipg_7/ffi_1/nand_6/w_0_0# gnd 0.10fF
C1553 ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_6/a 0.31fF
C1554 ffipg_4/ffi_1/nand_1/b ffipg_4/ffi_1/nand_3/b 0.32fF
C1555 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# 0.04fF
C1556 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C1557 nor_0/a nor_0/b 0.32fF
C1558 cla_2/p1 ffipg_3/k 0.05fF
C1559 clk ffipg_0/ffi_1/nand_3/a 0.13fF
C1560 gnd ffipg_0/ffi_0/nand_3/w_0_0# 0.11fF
C1561 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C1562 clk sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1563 sumffo_0/ffo_0/nand_7/a gnd 0.33fF
C1564 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C1565 ffipg_7/ffi_0/nand_6/a ffipg_7/ffi_0/qbar 0.00fF
C1566 ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_7/a 0.00fF
C1567 ffipg_4/ffi_1/inv_1/op ffipg_4/ffi_1/nand_4/w_0_0# 0.06fF
C1568 gnd ffipg_4/pggen_0/xor_0/w_n3_4# 0.12fF
C1569 gnd ffipg_1/ffi_0/inv_1/op 1.85fF
C1570 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C1571 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_1/b 0.04fF
C1572 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/nand_6/a 0.06fF
C1573 gnd ffipg_3/ffi_0/inv_0/op 0.27fF
C1574 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C1575 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C1576 inv_4/in cla_1/n 0.02fF
C1577 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C1578 ffipg_6/pggen_0/xor_0/a_10_10# ffipg_6/k 0.45fF
C1579 ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/nand_7/w_0_0# 0.06fF
C1580 ffipg_7/pggen_0/nand_0/w_0_0# gnd 0.10fF
C1581 clk sumffo_2/ffo_0/d 0.25fF
C1582 inv_0/op inv_0/in 0.04fF
C1583 sumffo_3/xor_0/w_n3_4# ffipg_3/k 0.06fF
C1584 sumffo_0/sbar sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C1585 sumffo_0/ffo_0/nand_6/w_0_0# z1o 0.06fF
C1586 ffipg_7/ffi_1/nand_3/a ffipg_7/ffi_1/nand_3/w_0_0# 0.06fF
C1587 ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/nand_1/w_0_0# 0.06fF
C1588 ffipg_7/ffi_1/nand_1/a gnd 0.44fF
C1589 ffipg_5/ffi_0/nand_6/a ffipg_5/ffi_0/qbar 0.00fF
C1590 gnd ffi_0/nand_6/w_0_0# 0.10fF
C1591 ffi_1/nand_2/w_0_0# ffi_1/nand_3/a 0.04fF
C1592 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b 0.32fF
C1593 nor_3/w_0_0# nor_4/b 0.03fF
C1594 gnd ffipg_4/ffi_1/nand_7/w_0_0# 0.10fF
C1595 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/a 0.06fF
C1596 gnd ffipg_4/pggen_0/xor_0/a_10_10# 0.93fF
C1597 gnd ffipg_3/ffi_1/inv_1/op 1.85fF
C1598 gnd ffipg_3/ffi_1/nand_2/w_0_0# 0.10fF
C1599 gnd cinin 0.44fF
C1600 clk ffipg_2/ffi_1/inv_0/op 0.32fF
C1601 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_6/a 0.13fF
C1602 clk ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C1603 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C1604 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_3/b 0.04fF
C1605 cla_2/p1 gnd 1.00fF
C1606 ffipg_7/ffi_0/inv_0/op ffipg_7/ffi_0/inv_0/w_0_6# 0.03fF
C1607 ffipg_7/ffi_0/nand_3/a ffipg_7/ffi_0/nand_3/w_0_0# 0.06fF
C1608 ffipg_4/ffi_1/nand_1/w_0_0# ffipg_4/ffi_1/nand_3/b 0.04fF
C1609 ffipg_2/ffi_1/nand_0/w_0_0# ffipg_2/ffi_1/nand_1/a 0.04fF
C1610 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/ffi_0/q 0.23fF
C1611 ffo_0/nand_0/w_0_0# ffo_0/nand_0/b 0.06fF
C1612 ffipg_4/ffi_0/inv_1/op ffipg_4/ffi_0/nand_1/b 0.45fF
C1613 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C1614 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_1/b 0.45fF
C1615 ffipg_7/ffi_1/nand_3/w_0_0# ffipg_7/ffi_1/nand_3/b 0.06fF
C1616 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C1617 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_7/a 0.04fF
C1618 ffipg_5/ffi_1/nand_6/a ffipg_5/ffi_1/qbar 0.00fF
C1619 ffipg_5/ffi_1/nand_4/w_0_0# ffipg_5/ffi_1/inv_1/op 0.06fF
C1620 gnd ffipg_5/ffi_0/nand_0/w_0_0# 0.10fF
C1621 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a 0.13fF
C1622 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/ffi_0/q 0.06fF
C1623 gnd ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C1624 gnd ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C1625 gnd inv_3/w_0_6# 0.17fF
C1626 ffipg_1/ffi_0/inv_0/op ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C1627 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/b 0.32fF
C1628 ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_0/nand_6/a 0.13fF
C1629 cla_2/nand_0/a_13_n26# gnd 0.01fF
C1630 gnd ffi_0/nand_6/a 0.33fF
C1631 clk ffipg_2/ffi_1/nand_3/a 0.13fF
C1632 ffo_0/inv_0/op ffo_0/nand_0/b 0.32fF
C1633 gnd sumffo_3/xor_0/w_n3_4# 0.12fF
C1634 ffipg_7/ffi_1/inv_1/op clk 0.07fF
C1635 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_3/w_0_0# 0.06fF
C1636 ffipg_6/ffi_1/q ffipg_6/k 0.46fF
C1637 ffipg_6/ffi_0/q ffipg_6/p 0.03fF
C1638 ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/pggen_0/xor_0/inv_1/op 0.08fF
C1639 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a 0.31fF
C1640 gnd ffo_0/nand_3/a 0.48fF
C1641 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C1642 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/nand_6/a 0.06fF
C1643 cla_0/nand_0/a_13_n26# gnd 0.00fF
C1644 clk y1in 1.36fF
C1645 sumffo_3/ffo_0/d sumffo_3/ffo_0/inv_0/op 0.04fF
C1646 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C1647 sumffo_0/ffo_0/nand_3/a gnd 0.33fF
C1648 cla_2/g1 cla_2/inv_0/op 0.35fF
C1649 ffipg_6/ffi_1/nand_3/a ffipg_6/ffi_1/nand_3/b 0.31fF
C1650 x2in ffipg_5/ffi_1/inv_1/op 0.01fF
C1651 ffi_0/inv_1/op ffi_0/inv_1/w_0_6# 0.04fF
C1652 gnd ffi_0/inv_0/op 0.27fF
C1653 ffipg_1/ffi_0/nand_3/w_0_0# ffipg_1/ffi_0/nand_3/b 0.06fF
C1654 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar 0.32fF
C1655 gnd ffipg_3/ffi_0/qbar 0.67fF
C1656 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C1657 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C1658 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C1659 cla_0/g0 cla_0/l 0.14fF
C1660 ffipg_6/ffi_1/nand_3/a gnd 0.33fF
C1661 ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_7/a 0.00fF
C1662 ffi_1/nand_1/b ffi_1/nand_7/a 0.13fF
C1663 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a 0.00fF
C1664 ffipg_2/ffi_0/q ffipg_2/ffi_1/q 0.73fF
C1665 ffipg_7/ffi_0/inv_1/op ffipg_7/ffi_0/nand_1/b 0.45fF
C1666 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C1667 clk ffi_0/nand_2/w_0_0# 0.06fF
C1668 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/a 0.31fF
C1669 ffipg_2/k sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C1670 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C1671 cla_0/l cla_2/p0 0.44fF
C1672 ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_6/w_0_0# 0.06fF
C1673 ffipg_6/pggen_0/xor_0/a_10_10# gnd 0.93fF
C1674 ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C1675 ffipg_2/ffi_0/nand_0/w_0_0# ffipg_2/ffi_0/nand_1/a 0.04fF
C1676 gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1677 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op 0.06fF
C1678 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/b 0.32fF
C1679 ffi_1/nand_7/a cinq 0.00fF
C1680 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/a 0.31fF
C1681 clk ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C1682 sumffo_3/ffo_0/nand_6/a sumffo_3/sbar 0.00fF
C1683 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C1684 nor_0/b ffi_0/nand_7/a 0.31fF
C1685 ffi_0/inv_1/op ffi_0/nand_3/b 0.33fF
C1686 clk ffi_0/nand_0/w_0_0# 0.06fF
C1687 gnd ffipg_3/ffi_0/nand_1/b 0.57fF
C1688 gnd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C1689 clk x1in 1.36fF
C1690 gnd sumffo_1/ffo_0/nand_2/w_0_0# 0.10fF
C1691 cla_0/l cla_1/n 0.13fF
C1692 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C1693 ffipg_6/ffi_0/inv_1/w_0_6# gnd 0.06fF
C1694 ffipg_4/pggen_0/xor_0/w_n3_4# ffipg_4/pggen_0/xor_0/inv_1/op 0.06fF
C1695 gnd ffipg_2/ffi_1/qbar 0.67fF
C1696 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1697 gnd ffipg_1/ffi_0/nand_1/a 0.44fF
C1698 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C1699 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C1700 ffipg_6/ffi_1/nand_3/a ffipg_6/ffi_1/nand_2/w_0_0# 0.04fF
C1701 ffipg_5/ffi_0/nand_3/a ffipg_5/ffi_0/nand_2/w_0_0# 0.04fF
C1702 clk ffi_0/inv_1/op 0.93fF
C1703 clk ffipg_2/ffi_1/inv_1/op 0.07fF
C1704 ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/nand_3/b 0.00fF
C1705 ffipg_7/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C1706 ffipg_7/ffi_0/nand_2/w_0_0# clk 0.06fF
C1707 ffipg_5/ffi_1/q ffipg_5/ffi_1/nand_6/a 0.31fF
C1708 ffipg_5/p ffipg_5/k 0.05fF
C1709 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_1/b 0.04fF
C1710 gnd ffo_0/nand_1/w_0_0# 0.10fF
C1711 gnd ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C1712 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C1713 gnd ffipg_4/ffi_1/nand_0/w_0_0# 0.10fF
C1714 ffipg_4/ffi_0/nand_4/w_0_0# ffipg_4/ffi_0/nand_3/b 0.06fF
C1715 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C1716 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_1/b 0.06fF
C1717 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C1718 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C1719 ffipg_5/pggen_0/xor_0/w_n3_4# ffipg_5/k 0.02fF
C1720 ffi_0/nand_3/a ffi_0/nand_2/w_0_0# 0.04fF
C1721 nor_4/b inv_9/in 0.16fF
C1722 ffipg_1/ffi_1/inv_0/op ffipg_1/ffi_1/inv_0/w_0_6# 0.03fF
C1723 gnd nor_2/b 0.32fF
C1724 clk sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C1725 gnd sumffo_2/ffo_0/nand_6/w_0_0# 0.10fF
C1726 ffipg_6/ffi_0/inv_0/w_0_6# gnd 0.06fF
C1727 ffipg_4/ffi_0/nand_4/w_0_0# ffipg_4/ffi_0/nand_6/a 0.04fF
C1728 y2in ffipg_5/ffi_0/inv_1/op 0.01fF
C1729 gnd ffipg_3/ffi_0/nand_1/w_0_0# 0.10fF
C1730 gnd ffi_1/nand_3/a 0.33fF
C1731 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a 0.00fF
C1732 gnd ffipg_0/ffi_1/nand_7/a 0.37fF
C1733 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1734 inv_1/op gnd 0.58fF
C1735 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/nand_0/b 0.06fF
C1736 cla_0/inv_0/in cla_0/inv_0/op 0.04fF
C1737 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C1738 ffipg_6/ffi_1/q gnd 2.24fF
C1739 gnd ffipg_4/ffi_1/nand_6/w_0_0# 0.10fF
C1740 ffipg_5/ffi_0/q ffipg_5/k 0.07fF
C1741 ffipg_2/ffi_1/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C1742 sumffo_2/xor_0/inv_1/op ffipg_2/k 0.22fF
C1743 ffi_0/q sumffo_2/xor_0/inv_0/op 0.06fF
C1744 gnd ffipg_1/ffi_0/qbar 0.67fF
C1745 sumffo_3/xor_0/a_10_10# ffipg_3/k 0.12fF
C1746 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C1747 gnd sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1748 ffipg_6/ffi_0/inv_1/op gnd 1.85fF
C1749 ffi_1/inv_1/op ffi_1/inv_1/w_0_6# 0.04fF
C1750 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_1/a 0.06fF
C1751 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_1/b 0.04fF
C1752 ffipg_0/ffi_1/nand_6/w_0_0# ffipg_0/ffi_1/nand_6/a 0.06fF
C1753 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C1754 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C1755 ffipg_6/ffi_1/nand_7/w_0_0# ffipg_6/ffi_1/qbar 0.06fF
C1756 gnd ffipg_4/ffi_0/nand_6/w_0_0# 0.10fF
C1757 clk ffipg_3/ffi_0/inv_1/op 0.07fF
C1758 gnd ffipg_0/ffi_0/nand_6/w_0_0# 0.10fF
C1759 gnd ffo_0/nand_7/w_0_0# 0.10fF
C1760 clk sumffo_1/ffo_0/nand_3/b 0.33fF
C1761 ffipg_7/ffi_0/qbar gnd 0.67fF
C1762 ffipg_6/ffi_0/nand_7/a gnd 0.37fF
C1763 gnd ffipg_3/ffi_1/nand_7/a 0.37fF
C1764 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a 0.31fF
C1765 clk ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C1766 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1767 ffo_0/nand_0/b ffo_0/nand_3/a 0.13fF
C1768 ffo_0/nand_1/a gnd 0.33fF
C1769 sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d 0.52fF
C1770 sumffo_0/ffo_0/nand_0/b clk 0.04fF
C1771 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C1772 ffipg_3/ffi_0/nand_2/w_0_0# y4in 0.06fF
C1773 ffi_0/q sumffo_3/xor_0/inv_1/op 0.04fF
C1774 ffipg_5/ffi_1/q ffipg_5/pggen_0/xor_0/inv_1/op 0.06fF
C1775 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C1776 y3in ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C1777 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C1778 cla_0/l inv_7/w_0_6# 0.06fF
C1779 gnd ffipg_1/ffi_0/nand_1/b 0.57fF
C1780 gnd ffipg_0/ffi_0/nand_3/a 0.33fF
C1781 sumffo_3/ffo_0/d gnd 0.41fF
C1782 clk sumffo_2/ffo_0/nand_3/b 0.33fF
C1783 cla_0/nor_1/w_0_0# gnd 0.31fF
C1784 gnd ffipg_4/ffi_0/nand_3/a 0.33fF
C1785 ffipg_4/ffi_1/q ffipg_4/pggen_0/xor_0/inv_0/op 0.27fF
C1786 ffipg_5/ffi_1/nand_4/w_0_0# ffipg_5/ffi_1/nand_6/a 0.04fF
C1787 ffipg_5/ffi_0/nand_7/w_0_0# ffipg_5/ffi_0/nand_7/a 0.06fF
C1788 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# 0.04fF
C1789 clk ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1790 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C1791 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a 0.13fF
C1792 ffi_0/nand_1/b ffi_0/nand_7/a 0.13fF
C1793 ffi_0/nand_5/w_0_0# ffi_0/inv_1/op 0.06fF
C1794 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/nand_6/a 0.06fF
C1795 gnd ffipg_1/ffi_1/inv_0/op 0.27fF
C1796 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q 0.27fF
C1797 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C1798 gnd sumffo_3/xor_0/a_10_10# 0.93fF
C1799 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b 0.13fF
C1800 cla_2/inv_0/in gnd 0.34fF
C1801 inv_0/op cla_0/g0 0.32fF
C1802 ffipg_7/ffi_1/nand_1/w_0_0# ffipg_7/ffi_1/nand_1/b 0.06fF
C1803 ffipg_7/ffi_1/nand_1/b gnd 0.57fF
C1804 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/nand_6/w_0_0# 0.06fF
C1805 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_7/a 0.13fF
C1806 gnd y3in 0.44fF
C1807 cla_1/inv_0/op cla_0/n 0.02fF
C1808 ffipg_0/ffi_0/nand_1/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C1809 gnd ffo_0/nand_6/w_0_0# 0.10fF
C1810 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_1/inv_1/op 0.75fF
C1811 inv_6/in nor_4/b 0.04fF
C1812 sumffo_0/sbar sumffo_0/ffo_0/nand_7/a 0.31fF
C1813 sumffo_0/ffo_0/nand_6/w_0_0# gnd 0.10fF
C1814 sumffo_0/ffo_0/nand_6/a z1o 0.31fF
C1815 cla_0/l cla_1/p0 0.09fF
C1816 ffipg_5/ffi_1/nand_7/w_0_0# ffipg_5/ffi_1/nand_7/a 0.06fF
C1817 gnd ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C1818 gnd x4in 0.44fF
C1819 ffipg_7/ffi_0/nand_6/w_0_0# ffipg_7/ffi_0/nand_6/a 0.06fF
C1820 sumffo_2/xor_0/inv_1/op ffi_0/q 0.04fF
C1821 nor_0/w_0_0# ffi_0/q 0.16fF
C1822 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/ffi_1/q 0.27fF
C1823 clk x2in 1.36fF
C1824 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C1825 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C1826 sumffo_1/ffo_0/nand_6/a clk 0.13fF
C1827 cla_2/nor_1/w_0_0# gnd 0.31fF
C1828 ffipg_7/ffi_1/nand_4/w_0_0# ffipg_7/ffi_1/nand_6/a 0.04fF
C1829 ffipg_7/ffi_0/inv_1/op gnd 1.85fF
C1830 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a 0.31fF
C1831 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/inv_1/op 0.06fF
C1832 nand_2/b inv_2/w_0_6# 0.03fF
C1833 clk ffipg_1/ffi_0/inv_1/op 0.07fF
C1834 gnd ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C1835 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C1836 gnd sumffo_1/ffo_0/nand_7/w_0_0# 0.10fF
C1837 sumffo_2/xor_0/w_n3_4# gnd 0.12fF
C1838 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C1839 ffipg_6/ffi_0/nand_3/a ffipg_6/ffi_0/nand_3/b 0.31fF
C1840 gnd ffipg_4/ffi_1/nand_6/a 0.37fF
C1841 ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/w_n3_4# 0.06fF
C1842 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C1843 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/inv_0/op 0.06fF
C1844 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/nand_3/b 0.06fF
C1845 gnd ffipg_5/p 0.35fF
C1846 gnd ffipg_2/ffi_0/nand_7/a 0.37fF
C1847 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C1848 cla_0/g0 cla_1/p0 0.38fF
C1849 ffipg_7/ffi_1/nand_1/a ffipg_7/ffi_1/nand_0/w_0_0# 0.04fF
C1850 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1851 ffipg_6/ffi_0/q ffipg_6/k 0.07fF
C1852 ffipg_4/ffi_1/nand_7/a ffipg_4/ffi_1/nand_5/w_0_0# 0.04fF
C1853 gnd ffipg_5/pggen_0/xor_0/w_n3_4# 0.12fF
C1854 clk ffipg_3/ffi_0/inv_0/op 0.32fF
C1855 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C1856 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/ffi_1/q 0.06fF
C1857 gnd sumffo_3/ffo_0/nand_0/b 0.53fF
C1858 cla_1/nor_1/w_0_0# gnd 0.31fF
C1859 cla_1/p0 cla_2/p0 0.24fF
C1860 ffipg_7/ffi_0/nand_1/w_0_0# ffipg_7/ffi_0/nand_1/a 0.06fF
C1861 ffipg_7/pggen_0/nor_0/w_0_0# ffipg_7/ffi_1/q 0.06fF
C1862 x1in ffipg_0/ffi_1/inv_1/op 0.01fF
C1863 gnd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C1864 gnd inv_0/in 0.30fF
C1865 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/d 0.06fF
C1866 ffipg_0/k gnd 0.68fF
C1867 ffipg_7/ffi_1/nand_1/a clk 0.13fF
C1868 ffipg_5/ffi_1/inv_0/op ffipg_5/ffi_1/inv_0/w_0_6# 0.03fF
C1869 gnd ffipg_5/ffi_1/nand_1/w_0_0# 0.10fF
C1870 ffipg_5/ffi_0/nand_5/w_0_0# ffipg_5/ffi_0/inv_1/op 0.06fF
C1871 ffi_1/inv_1/op ffi_1/nand_4/w_0_0# 0.06fF
C1872 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_1/b 0.45fF
C1873 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a 0.31fF
C1874 ffipg_1/ffi_1/nand_2/w_0_0# ffipg_1/ffi_1/nand_3/a 0.04fF
C1875 gnd ffipg_4/ffi_1/nand_5/w_0_0# 0.10fF
C1876 gnd ffipg_5/ffi_0/q 3.00fF
C1877 gnd ffi_1/nand_1/a 0.44fF
C1878 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a 0.00fF
C1879 ffo_0/nand_1/a ffo_0/nand_0/b 0.13fF
C1880 gnd sumffo_1/xor_0/inv_0/op 0.32fF
C1881 y2in ffipg_5/ffi_0/inv_0/w_0_6# 0.06fF
C1882 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/nand_6/a 0.04fF
C1883 ffipg_6/ffi_1/q ffipg_6/pggen_0/xor_0/inv_1/op 0.06fF
C1884 ffipg_4/ffi_0/q ffipg_4/pggen_0/xor_0/a_10_10# 0.12fF
C1885 clk ffipg_3/ffi_1/inv_1/op 0.07fF
C1886 clk ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C1887 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_1/b 0.04fF
C1888 ffi_0/q nor_0/b 0.32fF
C1889 clk cinin 1.36fF
C1890 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C1891 ffipg_6/ffi_0/nand_1/w_0_0# ffipg_6/ffi_0/nand_1/b 0.06fF
C1892 ffipg_5/ffi_1/q ffipg_5/pggen_0/nand_0/w_0_0# 0.06fF
C1893 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# 0.04fF
C1894 ffipg_1/ffi_0/nand_2/w_0_0# y2in 0.06fF
C1895 gnd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C1896 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_1/a 0.04fF
C1897 gnd sumffo_0/xor_0/a_10_10# 0.93fF
C1898 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1899 cla_1/inv_0/w_0_6# gnd 0.06fF
C1900 ffipg_6/ffi_1/nand_6/a ffipg_6/ffi_1/nand_4/w_0_0# 0.04fF
C1901 ffipg_6/ffi_0/inv_1/op ffipg_6/ffi_0/nand_6/a 0.13fF
C1902 ffipg_5/ffi_1/nand_3/w_0_0# ffipg_5/ffi_1/nand_3/b 0.06fF
C1903 gnd ffipg_5/ffi_1/nand_3/b 0.74fF
C1904 clk ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C1905 ffipg_7/ffi_1/nand_3/b ffipg_7/ffi_1/nand_1/b 0.32fF
C1906 clk ffipg_5/ffi_0/nand_0/w_0_0# 0.06fF
C1907 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_0/q 0.06fF
C1908 gnd inv_4/in 0.33fF
C1909 gnd z3o 0.80fF
C1910 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b 0.32fF
C1911 cla_0/nor_0/w_0_0# gnd 0.31fF
C1912 ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_6/w_0_0# 0.06fF
C1913 gnd ffipg_5/ffi_1/nand_2/w_0_0# 0.10fF
C1914 gnd ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C1915 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C1916 sumffo_1/ffo_0/inv_0/op gnd 0.27fF
C1917 ffipg_7/ffi_1/nand_2/w_0_0# x4in 0.06fF
C1918 ffipg_7/ffi_0/nand_4/w_0_0# ffipg_7/ffi_0/nand_6/a 0.04fF
C1919 ffipg_6/ffi_0/q ffipg_6/g 0.13fF
C1920 ffi_0/q sumffo_1/xor_0/a_10_10# 0.04fF
C1921 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_3/b 0.00fF
C1922 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/nand_7/a 0.06fF
C1923 ffipg_7/ffi_0/nand_7/w_0_0# ffipg_7/ffi_0/nand_7/a 0.06fF
C1924 ffipg_6/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C1925 gnd ffipg_4/ffi_1/inv_1/w_0_6# 0.06fF
C1926 ffipg_4/ffi_1/nand_1/w_0_0# ffipg_4/ffi_1/nand_1/b 0.06fF
C1927 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_1/a 0.06fF
C1928 gnd nor_4/a 0.40fF
C1929 cla_1/nand_0/a_13_n26# gnd 0.01fF
C1930 gnd ffi_1/inv_0/w_0_6# 0.06fF
C1931 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C1932 gnd sumffo_2/ffo_0/nand_0/b 0.63fF
C1933 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/inv_1/w_0_6# 0.04fF
C1934 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a 0.31fF
C1935 clk ffi_0/inv_0/op 0.32fF
C1936 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C1937 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/inv_1/op 0.33fF
C1938 ffipg_7/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1939 y1in ffipg_4/ffi_0/inv_0/w_0_6# 0.06fF
C1940 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_3/b 0.00fF
C1941 gnd ffipg_3/ffi_0/nand_4/w_0_0# 0.10fF
C1942 ffipg_3/ffi_1/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C1943 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_1/op 0.08fF
C1944 y1in ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1945 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_6/a 0.04fF
C1946 ffipg_3/k inv_4/op 0.09fF
C1947 gnd sumffo_2/ffo_0/nand_6/a 0.33fF
C1948 ffipg_6/ffi_1/nand_3/a clk 0.13fF
C1949 ffipg_7/ffi_1/inv_0/w_0_6# x4in 0.06fF
C1950 ffo_0/nand_7/w_0_0# couto 0.04fF
C1951 ffipg_6/ffi_0/q gnd 3.00fF
C1952 gnd ffipg_4/ffi_1/nand_4/w_0_0# 0.10fF
C1953 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b 0.32fF
C1954 gnd ffipg_1/ffi_1/nand_7/w_0_0# 0.10fF
C1955 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C1956 ffipg_6/ffi_1/inv_1/op x3in 0.01fF
C1957 gnd ffi_1/qbar 0.62fF
C1958 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_7/a 0.04fF
C1959 y1in ffipg_0/ffi_0/inv_1/op 0.01fF
C1960 ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_3/b 0.31fF
C1961 gnd sumffo_3/ffo_0/nand_0/w_0_0# 0.10fF
C1962 ffipg_7/ffi_1/nand_6/w_0_0# ffipg_7/ffi_1/qbar 0.04fF
C1963 ffipg_7/ffi_1/nand_1/b ffipg_7/ffi_1/nand_7/a 0.13fF
C1964 y1in ffipg_4/ffi_0/inv_1/op 0.01fF
C1965 gnd ffipg_4/ffi_0/nand_4/w_0_0# 0.10fF
C1966 ffipg_5/ffi_1/nand_3/a ffipg_5/ffi_1/nand_3/b 0.31fF
C1967 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_0/q 0.20fF
C1968 ffi_1/nand_3/w_0_0# ffi_1/nand_1/b 0.04fF
C1969 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a 0.13fF
C1970 cla_2/l cla_0/n 0.32fF
C1971 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C1972 ffipg_6/ffi_1/nand_1/b ffipg_6/ffi_1/nand_3/b 0.32fF
C1973 ffi_0/nand_4/w_0_0# ffi_0/inv_1/op 0.06fF
C1974 gnd ffo_0/nand_7/a 0.33fF
C1975 ffipg_7/k ffipg_7/pggen_0/nor_0/a_13_6# 0.01fF
C1976 ffipg_6/ffi_1/nand_1/b gnd 0.57fF
C1977 ffipg_6/ffi_0/inv_1/w_0_6# clk 0.06fF
C1978 ffipg_7/pggen_0/xor_0/inv_1/w_0_6# ffipg_7/ffi_0/q 0.23fF
C1979 cla_0/l ffipg_3/k 0.10fF
C1980 ffipg_5/ffi_1/nand_2/w_0_0# ffipg_5/ffi_1/nand_3/a 0.04fF
C1981 ffipg_5/ffi_1/nand_1/a ffipg_5/ffi_1/nand_1/b 0.31fF
C1982 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/inv_1/w_0_6# 0.04fF
C1983 ffi_1/nand_1/b ffi_1/inv_1/op 0.45fF
C1984 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C1985 clk ffipg_1/ffi_0/nand_1/a 0.13fF
C1986 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C1987 gnd ffipg_0/ffi_1/nand_6/w_0_0# 0.10fF
C1988 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C1989 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C1990 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_1/op 0.52fF
C1991 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a 0.00fF
C1992 ffipg_7/ffi_1/nand_6/a gnd 0.37fF
C1993 ffipg_7/ffi_0/q ffipg_7/ffi_0/nand_7/w_0_0# 0.04fF
C1994 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a 0.00fF
C1995 inv_5/in nor_3/b 0.04fF
C1996 gnd inv_4/op 0.58fF
C1997 cla_0/l inv_7/in 0.13fF
C1998 ffipg_6/ffi_1/nand_6/w_0_0# gnd 0.10fF
C1999 gnd ffipg_2/ffi_0/nand_4/w_0_0# 0.10fF
C2000 gnd inv_5/in 0.49fF
C2001 nand_2/b cla_0/n 0.00fF
C2002 gnd ffipg_5/ffi_0/nand_7/w_0_0# 0.10fF
C2003 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C2004 ffipg_2/ffi_0/q ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C2005 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C2006 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C2007 ffo_0/nand_6/w_0_0# couto 0.06fF
C2008 ffipg_7/k ffipg_7/ffi_1/q 0.46fF
C2009 ffipg_7/pggen_0/xor_0/inv_0/op ffipg_7/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C2010 clk ffipg_4/ffi_1/nand_0/w_0_0# 0.06fF
C2011 ffi_0/q sumffo_1/ffo_0/d 0.27fF
C2012 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_3/a 0.04fF
C2013 ffipg_6/ffi_1/inv_0/op ffipg_6/ffi_1/inv_0/w_0_6# 0.03fF
C2014 ffipg_6/p ffipg_6/k 0.05fF
C2015 gnd ffipg_5/ffi_1/nand_7/w_0_0# 0.10fF
C2016 ffipg_5/ffi_1/nand_3/b ffipg_5/ffi_1/inv_1/op 0.33fF
C2017 ffipg_5/g ffipg_5/ffi_0/q 0.13fF
C2018 gnd ffipg_3/ffi_1/nand_6/w_0_0# 0.10fF
C2019 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a 0.31fF
C2020 gnd ffipg_3/ffi_1/inv_0/op 0.27fF
C2021 clk ffi_1/nand_3/a 0.13fF
C2022 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_7/a 0.04fF
C2023 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C2024 ffo_0/nand_2/w_0_0# ffo_0/d 0.06fF
C2025 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C2026 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C2027 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C2028 ffipg_7/ffi_0/nand_3/a ffipg_7/ffi_0/nand_2/w_0_0# 0.04fF
C2029 gnd ffo_0/nand_6/a 0.33fF
C2030 ffipg_7/ffi_0/nand_6/w_0_0# gnd 0.10fF
C2031 ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/nand_1/w_0_0# 0.06fF
C2032 ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C2033 x1in ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C2034 ffipg_7/pggen_0/nor_0/w_0_0# ffipg_7/k 0.21fF
C2035 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C2036 ffipg_0/k ffipg_0/ffi_1/q 0.46fF
C2037 cla_2/p0 ffipg_3/k 0.06fF
C2038 gnd ffi_1/nand_3/b 0.74fF
C2039 gnd ffipg_1/ffi_0/nand_4/w_0_0# 0.10fF
C2040 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C2041 gnd ffipg_0/ffi_1/nand_2/w_0_0# 0.10fF
C2042 cla_2/n nor_3/b 0.41fF
C2043 ffo_0/nand_5/w_0_0# ffo_0/nand_7/a 0.04fF
C2044 clk sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C2045 sumffo_0/ffo_0/nand_6/a gnd 0.33fF
C2046 cla_0/l gnd 3.05fF
C2047 ffipg_6/ffi_0/inv_1/op clk 0.07fF
C2048 ffipg_6/ffi_0/nand_4/w_0_0# ffipg_6/ffi_0/nand_3/b 0.06fF
C2049 x1in ffipg_4/ffi_1/inv_0/w_0_6# 0.06fF
C2050 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/nand_6/a 0.06fF
C2051 ffi_1/inv_1/op ffi_1/nand_6/a 0.13fF
C2052 gnd ffipg_4/ffi_1/inv_1/op 1.85fF
C2053 gnd cla_2/n 0.60fF
C2054 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C2055 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_1/op 0.06fF
C2056 ffipg_4/ffi_0/q ffipg_4/ffi_0/nand_6/w_0_0# 0.06fF
C2057 gnd ffipg_4/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C2058 ffipg_4/ffi_1/q ffipg_4/pggen_0/nand_0/w_0_0# 0.06fF
C2059 gnd ffipg_3/ffi_1/nand_1/b 0.57fF
C2060 ffi_0/nand_7/w_0_0# nor_0/b 0.06fF
C2061 ffi_0/nand_1/b ffi_0/inv_1/op 0.45fF
C2062 ffi_1/nand_1/a ffi_1/nand_0/w_0_0# 0.04fF
C2063 cla_1/inv_0/in cla_1/inv_0/w_0_6# 0.06fF
C2064 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C2065 clk sumffo_3/ffo_0/d 0.04fF
C2066 clk ffipg_4/ffi_0/nand_3/a 0.13fF
C2067 clk ffipg_0/ffi_0/nand_3/a 0.13fF
C2068 ffi_0/q sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C2069 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/sbar 0.04fF
C2070 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a 0.13fF
C2071 x1in ffipg_4/ffi_1/nand_2/w_0_0# 0.06fF
C2072 x1in ffipg_4/ffi_1/inv_0/op 0.04fF
C2073 gnd ffipg_2/ffi_1/nand_3/w_0_0# 0.11fF
C2074 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/inv_1/w_0_6# 0.04fF
C2075 sumffo_1/sbar z2o 0.32fF
C2076 gnd sumffo_1/ffo_0/nand_4/w_0_0# 0.10fF
C2077 cla_0/g0 gnd 1.11fF
C2078 ffipg_7/ffi_1/q ffipg_7/pggen_0/xor_0/w_n3_4# 0.06fF
C2079 ffipg_7/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C2080 ffipg_6/ffi_1/inv_0/w_0_6# x3in 0.06fF
C2081 ffipg_6/pggen_0/xor_0/inv_0/op ffipg_6/pggen_0/xor_0/w_n3_4# 0.06fF
C2082 ffipg_6/pggen_0/xor_0/inv_1/w_0_6# ffipg_6/pggen_0/xor_0/inv_1/op 0.03fF
C2083 gnd ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C2084 clk ffipg_1/ffi_1/inv_0/op 0.32fF
C2085 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b 0.13fF
C2086 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C2087 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/ffo_0/nand_7/a 0.06fF
C2088 sumffo_2/sbar z3o 0.32fF
C2089 cla_2/p0 gnd 1.06fF
C2090 clk y3in 1.36fF
C2091 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C2092 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C2093 gnd ffipg_4/k 0.27fF
C2094 gnd ffipg_5/ffi_0/nand_3/b 0.74fF
C2095 ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C2096 gnd ffipg_0/ffi_0/nand_0/w_0_0# 0.10fF
C2097 sumffo_3/sbar sumffo_3/ffo_0/nand_7/a 0.31fF
C2098 ffipg_7/ffi_1/inv_1/w_0_6# gnd 0.06fF
C2099 ffipg_6/ffi_1/nand_4/w_0_0# ffipg_6/ffi_1/nand_3/b 0.06fF
C2100 ffipg_6/ffi_0/nand_2/w_0_0# gnd 0.10fF
C2101 ffipg_4/ffi_1/q ffipg_4/ffi_1/qbar 0.32fF
C2102 y1in ffipg_4/ffi_0/nand_2/w_0_0# 0.06fF
C2103 x2in ffipg_5/ffi_1/inv_0/op 0.04fF
C2104 ffipg_5/ffi_0/nand_5/w_0_0# ffipg_5/ffi_0/nand_1/b 0.06fF
C2105 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C2106 gnd ffipg_2/ffi_0/qbar 0.67fF
C2107 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C2108 gnd ffipg_0/ffi_1/nand_0/w_0_0# 0.10fF
C2109 gnd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C2110 gnd cla_1/n 0.51fF
C2111 clk x4in 1.36fF
C2112 ffipg_6/ffi_1/nand_4/w_0_0# gnd 0.10fF
C2113 ffipg_4/ffi_0/nand_1/a ffipg_4/ffi_0/nand_3/b 0.00fF
C2114 ffipg_4/ffi_0/nand_1/w_0_0# ffipg_4/ffi_0/nand_1/b 0.06fF
C2115 inv_1/op sumffo_2/xor_0/inv_0/op 0.27fF
C2116 sumffo_3/xor_0/inv_0/w_0_6# inv_4/op 0.06fF
C2117 ffipg_7/ffi_0/nand_3/b ffipg_7/ffi_0/nand_1/w_0_0# 0.04fF
C2118 ffipg_6/ffi_0/q ffipg_6/pggen_0/xor_0/inv_1/op 0.22fF
C2119 ffipg_6/pggen_0/xor_0/inv_0/w_0_6# ffipg_6/pggen_0/xor_0/inv_0/op 0.03fF
C2120 p1 ffipg_4/k 0.05fF
C2121 ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C2122 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C2123 gnd ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C2124 gnd ffo_0/nand_2/w_0_0# 0.10fF
C2125 ffipg_7/ffi_0/inv_1/op clk 0.07fF
C2126 ffipg_7/ffi_0/nand_4/w_0_0# gnd 0.10fF
C2127 ffipg_6/ffi_1/q ffipg_6/ffi_1/nand_7/w_0_0# 0.04fF
C2128 ffipg_6/ffi_0/q ffipg_6/ffi_0/nand_6/a 0.31fF
C2129 ffipg_6/p gnd 0.35fF
C2130 gnd ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C2131 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C2132 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/b 0.32fF
C2133 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C2134 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/w_0_0# 0.06fF
C2135 cla_2/g1 cla_2/p1 0.00fF
C2136 ffipg_5/ffi_0/q ffipg_5/ffi_0/nand_6/a 0.31fF
C2137 gnd ffipg_5/ffi_0/inv_0/op 0.27fF
C2138 ffipg_5/ffi_0/nand_1/a ffipg_5/ffi_0/nand_1/b 0.31fF
C2139 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_7/a 0.04fF
C2140 ffipg_1/k ffipg_1/ffi_1/q 0.46fF
C2141 gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C2142 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C2143 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# 0.04fF
C2144 ffipg_6/ffi_1/inv_0/op x3in 0.04fF
C2145 gnd ffipg_5/ffi_0/nand_0/a_13_n26# 0.01fF
C2146 gnd ffipg_4/ffi_0/inv_0/op 0.27fF
C2147 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C2148 y2in ffipg_1/ffi_0/inv_1/op 0.01fF
C2149 sumffo_0/xor_0/inv_0/op gnd 0.32fF
C2150 nand_2/b ffipg_2/k 0.06fF
C2151 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# 0.04fF
C2152 clk sumffo_3/ffo_0/nand_0/b 0.04fF
C2153 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C2154 inv_7/w_0_6# inv_7/in 0.10fF
C2155 ffipg_7/ffi_0/inv_0/w_0_6# y4in 0.06fF
C2156 ffi_0/q inv_2/w_0_6# 0.06fF
C2157 ffipg_6/ffi_0/nand_1/w_0_0# gnd 0.10fF
C2158 ffipg_3/k ffipg_3/ffi_1/q 0.46fF
C2159 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C2160 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C2161 gnd ffipg_2/ffi_1/nand_2/w_0_0# 0.10fF
C2162 ffipg_1/ffi_0/nand_2/w_0_0# ffipg_1/ffi_0/nand_3/a 0.04fF
C2163 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C2164 gnd sumffo_1/ffo_0/nand_0/b 0.62fF
C2165 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C2166 ffipg_6/ffi_0/nand_6/w_0_0# gnd 0.10fF
C2167 ffipg_4/ffi_0/nand_3/w_0_0# ffipg_4/ffi_0/nand_1/b 0.04fF
C2168 ffi_1/qbar ffi_1/nand_7/w_0_0# 0.06fF
C2169 ffi_1/nand_6/w_0_0# cinq 0.06fF
C2170 ffipg_7/ffi_1/q ffipg_7/ffi_0/q 0.73fF
C2171 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C2172 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a 0.13fF
C2173 ffi_0/nand_6/a nor_0/b 0.00fF
C2174 gnd ffipg_3/ffi_0/nand_3/b 0.74fF
C2175 clk ffi_1/nand_1/a 0.13fF
C2176 gnd ffo_0/inv_1/w_0_6# 0.06fF
C2177 sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# 0.02fF
C2178 inv_0/op gnd 0.27fF
C2179 gnd ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C2180 cla_0/l ffipg_2/ffi_0/q 0.13fF
C2181 gnd ffipg_1/ffi_1/nand_5/w_0_0# 0.10fF
C2182 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C2183 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C2184 ffo_0/nand_3/w_0_0# ffo_0/nand_3/b 0.06fF
C2185 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C2186 ffipg_7/ffi_1/nand_7/w_0_0# gnd 0.10fF
C2187 cla_2/l inv_5/w_0_6# 0.08fF
C2188 ffipg_5/pggen_0/xor_0/w_n3_4# ffipg_5/pggen_0/xor_0/a_10_10# 0.16fF
C2189 ffo_0/nand_7/a couto 0.00fF
C2190 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C2191 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_1/op 0.52fF
C2192 gnd inv_7/w_0_6# 0.15fF
C2193 ffipg_6/ffi_1/inv_1/w_0_6# gnd 0.06fF
C2194 y3in ffipg_2/ffi_0/inv_1/op 0.01fF
C2195 ffipg_0/ffi_1/nand_0/w_0_0# ffipg_0/ffi_1/inv_0/op 0.06fF
C2196 gnd ffipg_4/ffi_0/nand_3/b 0.74fF
C2197 gnd ffipg_5/ffi_1/nand_0/w_0_0# 0.10fF
C2198 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C2199 ffipg_1/ffi_0/nand_6/w_0_0# ffipg_1/ffi_0/qbar 0.04fF
C2200 gnd ffipg_0/ffi_0/nand_4/w_0_0# 0.10fF
C2201 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C2202 sumffo_2/xor_0/inv_1/op inv_1/op 0.06fF
C2203 gnd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C2204 cla_0/l cla_1/inv_0/in 0.23fF
C2205 ffipg_7/pggen_0/nor_0/w_0_0# ffipg_7/ffi_0/q 0.06fF
C2206 ffipg_6/ffi_0/nand_1/b gnd 0.57fF
C2207 ffipg_3/ffi_0/inv_0/op ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C2208 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_0/q 0.12fF
C2209 ffi_1/nand_6/w_0_0# ffi_1/nand_6/a 0.06fF
C2210 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C2211 ffipg_5/pggen_0/xor_0/inv_1/op ffipg_5/pggen_0/xor_0/w_n3_4# 0.06fF
C2212 ffi_0/nand_4/w_0_0# ffi_0/nand_6/a 0.04fF
C2213 cla_0/inv_0/op nand_2/b 0.09fF
C2214 gnd ffipg_4/ffi_0/nand_6/a 0.37fF
C2215 ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/a_10_10# 0.12fF
C2216 gnd ffipg_3/ffi_1/q 2.24fF
C2217 gnd ffipg_0/ffi_0/nand_6/a 0.37fF
C2218 clk ffipg_5/ffi_1/nand_2/w_0_0# 0.06fF
C2219 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a 0.31fF
C2220 clk ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C2221 gnd ffipg_0/ffi_1/nand_6/a 0.37fF
C2222 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C2223 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C2224 ffipg_5/ffi_0/nand_3/w_0_0# ffipg_5/ffi_0/nand_3/b 0.06fF
C2225 clk nor_4/a 0.03fF
C2226 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C2227 gnd ffipg_4/ffi_1/nand_0/a_13_n26# 0.01fF
C2228 clk ffipg_4/ffi_1/inv_1/w_0_6# 0.06fF
C2229 ffipg_5/ffi_0/q ffipg_5/pggen_0/xor_0/inv_1/op 0.22fF
C2230 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a 0.31fF
C2231 ffipg_2/k cla_0/n 0.06fF
C2232 gnd ffipg_4/ffi_1/nand_1/a 0.45fF
C2233 gnd ffipg_5/ffi_0/nand_7/a 0.37fF
C2234 gnd ffipg_3/ffi_0/nand_1/a 0.45fF
C2235 cla_2/p0 ffipg_2/ffi_0/q 0.03fF
C2236 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a 0.13fF
C2237 gnd ffipg_0/ffi_1/nand_1/w_0_0# 0.10fF
C2238 ffo_0/nand_6/a couto 0.31fF
C2239 gnd sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C2240 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_0/op 0.06fF
C2241 clk sumffo_2/ffo_0/nand_0/b 0.04fF
C2242 z1o gnd 0.80fF
C2243 cla_1/p0 gnd 1.06fF
C2244 ffipg_4/pggen_0/xor_0/w_n3_4# ffipg_4/pggen_0/xor_0/inv_0/op 0.06fF
C2245 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C2246 ffi_0/q nand_2/b 0.04fF
C2247 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C2248 ffipg_7/k ffipg_7/pggen_0/xor_0/w_n3_4# 0.02fF
C2249 ffipg_1/k nor_0/a 0.06fF
C2250 ffipg_4/pggen_0/xor_0/inv_1/op ffipg_4/k 0.52fF
C2251 ffipg_5/ffi_1/nand_5/w_0_0# ffipg_5/ffi_1/nand_1/b 0.06fF
C2252 gnd ffipg_5/ffi_1/nand_7/a 0.37fF
C2253 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/qbar 0.04fF
C2254 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C2255 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C2256 gnd z4o 0.80fF
C2257 sumffo_2/ffo_0/nand_0/w_0_0# gnd 0.10fF
C2258 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C2259 cla_1/inv_0/in cla_2/p0 0.02fF
C2260 gnd ffipg_0/ffi_0/nand_1/a 0.44fF
C2261 ffipg_7/ffi_0/nand_6/a gnd 0.37fF
C2262 ffipg_6/ffi_1/nand_6/a gnd 0.37fF
C2263 ffipg_2/ffi_1/nand_0/w_0_0# ffipg_2/ffi_1/inv_0/op 0.06fF
C2264 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar 0.32fF
C2265 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C2266 ffipg_0/k ffipg_0/ffi_0/q 0.07fF
C2267 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/pggen_0/xor_0/w_n3_4# 0.06fF
C2268 ffipg_2/ffi_0/nand_0/w_0_0# ffipg_2/ffi_0/inv_0/op 0.06fF
C2269 cla_2/p1 ffipg_3/ffi_0/q 0.03fF
C2270 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a 0.13fF
C2271 gnd ffipg_1/ffi_0/nand_3/b 0.74fF
C2272 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C2273 cla_0/n nor_1/w_0_0# 0.06fF
C2274 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C2275 gnd sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C2276 sumffo_1/ffo_0/nand_1/w_0_0# gnd 0.10fF
C2277 nand_2/b inv_3/in 0.13fF
C2278 ffipg_6/ffi_1/nand_0/w_0_0# gnd 0.10fF
C2279 ffipg_6/ffi_0/nand_3/w_0_0# ffipg_6/ffi_0/nand_1/b 0.04fF
C2280 ffi_1/nand_4/w_0_0# ffi_1/nand_6/a 0.04fF
C2281 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C2282 gnd sumffo_2/xor_0/a_10_10# 0.93fF
C2283 ffipg_6/ffi_1/nand_7/a gnd 0.37fF
C2284 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C2285 ffipg_6/pggen_0/xor_0/w_n3_4# ffipg_6/pggen_0/xor_0/a_10_10# 0.16fF
C2286 ffipg_5/pggen_0/xor_0/inv_0/op ffipg_5/ffi_0/q 0.20fF
C2287 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a 0.13fF
C2288 ffipg_1/ffi_0/q ffipg_1/ffi_1/q 0.73fF
C2289 ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C2290 nand_2/b ffipg_1/k 0.15fF
C2291 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_3/a 0.04fF
C2292 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C2293 ffipg_7/ffi_0/nand_1/b gnd 0.57fF
C2294 ffipg_7/ffi_1/q ffipg_7/p 0.22fF
C2295 ffipg_6/ffi_0/nand_0/w_0_0# gnd 0.10fF
C2296 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C2297 cla_0/n inv_5/w_0_6# 0.06fF
C2298 cla_1/l nand_2/b 0.31fF
C2299 ffi_0/q sumffo_1/xor_0/a_38_n43# 0.01fF
C2300 inv_2/in nor_1/b 0.04fF
C2301 ffo_0/nand_0/b ffo_0/inv_1/w_0_6# 0.03fF
C2302 gnd sumffo_1/ffo_0/nand_7/a 0.33fF
C2303 sumffo_0/ffo_0/nand_6/a sumffo_0/sbar 0.00fF
C2304 cla_0/inv_0/w_0_6# gnd 0.06fF
C2305 ffipg_7/ffi_1/nand_5/w_0_0# ffipg_7/ffi_1/inv_1/op 0.06fF
C2306 ffipg_6/ffi_1/nand_1/w_0_0# ffipg_6/ffi_1/nand_1/b 0.06fF
C2307 gnd ffipg_4/ffi_1/nand_3/w_0_0# 0.11fF
C2308 ffipg_7/ffi_1/nand_4/w_0_0# gnd 0.10fF
C2309 y2in ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C2310 cla_0/n inv_1/in 0.02fF
C2311 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C2312 ffipg_7/pggen_0/nor_0/w_0_0# ffipg_7/p 0.05fF
C2313 ffipg_5/pggen_0/nor_0/w_0_0# ffipg_5/ffi_1/q 0.06fF
C2314 gnd ffipg_5/k 0.27fF
C2315 clk ffipg_3/ffi_1/inv_0/op 0.32fF
C2316 gnd ffi_1/nand_2/w_0_0# 0.10fF
C2317 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C2318 gnd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C2319 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C2320 ffipg_4/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2321 ffipg_4/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2322 ffipg_4/ffi_1/nand_7/a Gnd 0.30fF
C2323 ffipg_4/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2324 ffipg_4/ffi_1/qbar Gnd 0.42fF
C2325 ffipg_4/ffi_1/nand_6/a Gnd 0.30fF
C2326 ffipg_4/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2327 ffipg_4/ffi_1/inv_1/op Gnd 0.89fF
C2328 ffipg_4/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2329 ffipg_4/ffi_1/nand_3/b Gnd 0.43fF
C2330 ffipg_4/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2331 ffipg_4/ffi_1/nand_3/a Gnd 0.30fF
C2332 ffipg_4/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2333 ffipg_4/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2334 ffipg_4/ffi_1/inv_0/op Gnd 0.26fF
C2335 ffipg_4/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2336 ffipg_4/ffi_1/nand_1/a Gnd 0.30fF
C2337 ffipg_4/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2338 ffipg_4/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2339 ffipg_4/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2340 ffipg_4/ffi_0/nand_7/a Gnd 0.30fF
C2341 ffipg_4/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2342 ffipg_4/ffi_0/qbar Gnd 0.42fF
C2343 ffipg_4/ffi_0/nand_6/a Gnd 0.30fF
C2344 ffipg_4/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2345 ffipg_4/ffi_0/inv_1/op Gnd 0.89fF
C2346 ffipg_4/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2347 ffipg_4/ffi_0/nand_3/b Gnd 0.43fF
C2348 ffipg_4/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2349 ffipg_4/ffi_0/nand_3/a Gnd 0.30fF
C2350 ffipg_4/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2351 ffipg_4/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2352 ffipg_4/ffi_0/inv_0/op Gnd 0.26fF
C2353 ffipg_4/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2354 ffipg_4/ffi_0/nand_1/a Gnd 0.30fF
C2355 ffipg_4/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2356 p1 Gnd 0.46fF
C2357 ffipg_4/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2358 ffipg_4/k Gnd 1.09fF
C2359 ffipg_4/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2360 ffipg_4/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2361 ffipg_4/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2362 ffipg_4/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2363 ffipg_4/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2364 ffipg_4/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2365 ffipg_4/g Gnd 0.13fF
C2366 ffipg_4/ffi_0/q Gnd 2.68fF
C2367 ffipg_4/ffi_1/q Gnd 2.93fF
C2368 ffipg_4/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2369 ffipg_5/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2370 ffipg_5/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2371 ffipg_5/ffi_1/nand_7/a Gnd 0.30fF
C2372 ffipg_5/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2373 ffipg_5/ffi_1/qbar Gnd 0.42fF
C2374 ffipg_5/ffi_1/nand_6/a Gnd 0.30fF
C2375 ffipg_5/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2376 ffipg_5/ffi_1/inv_1/op Gnd 0.89fF
C2377 ffipg_5/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2378 ffipg_5/ffi_1/nand_3/b Gnd 0.43fF
C2379 ffipg_5/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2380 ffipg_5/ffi_1/nand_3/a Gnd 0.30fF
C2381 ffipg_5/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2382 ffipg_5/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2383 ffipg_5/ffi_1/inv_0/op Gnd 0.26fF
C2384 ffipg_5/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2385 ffipg_5/ffi_1/nand_1/a Gnd 0.30fF
C2386 ffipg_5/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2387 ffipg_5/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2388 ffipg_5/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2389 ffipg_5/ffi_0/nand_7/a Gnd 0.30fF
C2390 ffipg_5/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2391 ffipg_5/ffi_0/qbar Gnd 0.42fF
C2392 ffipg_5/ffi_0/nand_6/a Gnd 0.30fF
C2393 ffipg_5/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2394 ffipg_5/ffi_0/inv_1/op Gnd 0.89fF
C2395 ffipg_5/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2396 ffipg_5/ffi_0/nand_3/b Gnd 0.43fF
C2397 ffipg_5/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2398 ffipg_5/ffi_0/nand_3/a Gnd 0.30fF
C2399 ffipg_5/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2400 ffipg_5/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2401 ffipg_5/ffi_0/inv_0/op Gnd 0.26fF
C2402 ffipg_5/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2403 ffipg_5/ffi_0/nand_1/a Gnd 0.30fF
C2404 ffipg_5/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2405 ffipg_5/p Gnd 0.46fF
C2406 ffipg_5/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2407 ffipg_5/k Gnd 1.09fF
C2408 ffipg_5/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2409 ffipg_5/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2410 ffipg_5/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2411 ffipg_5/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2412 ffipg_5/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2413 ffipg_5/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2414 ffipg_5/g Gnd 0.16fF
C2415 ffipg_5/ffi_0/q Gnd 2.68fF
C2416 ffipg_5/ffi_1/q Gnd 2.93fF
C2417 ffipg_5/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2418 ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2419 ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2420 ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C2421 ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2422 ffipg_3/ffi_1/qbar Gnd 0.42fF
C2423 ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C2424 ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2425 ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C2426 ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2427 ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C2428 ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2429 ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C2430 ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2431 x4in Gnd 1.03fF
C2432 ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2433 ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C2434 ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2435 ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C2436 ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2437 ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2438 ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2439 ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C2440 ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2441 ffipg_3/ffi_0/qbar Gnd 0.42fF
C2442 ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C2443 ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2444 ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C2445 ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2446 ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C2447 ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2448 ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C2449 ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2450 y4in Gnd 1.03fF
C2451 ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2452 ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C2453 ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2454 ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C2455 ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2456 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2457 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2458 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2459 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2460 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2461 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2462 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2463 ffipg_3/ffi_0/q Gnd 2.68fF
C2464 ffipg_3/ffi_1/q Gnd 2.93fF
C2465 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2466 ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2467 ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2468 ffi_0/nand_7/a Gnd 0.30fF
C2469 ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2470 nor_0/b Gnd 1.26fF
C2471 ffi_0/nand_6/a Gnd 0.30fF
C2472 ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2473 ffi_0/inv_1/op Gnd 0.89fF
C2474 ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2475 ffi_0/nand_3/b Gnd 0.43fF
C2476 ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2477 ffi_0/nand_3/a Gnd 0.30fF
C2478 ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2479 cinin Gnd 1.02fF
C2480 ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2481 ffi_0/inv_0/op Gnd 0.26fF
C2482 ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2483 ffi_0/nand_1/a Gnd 0.30fF
C2484 ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2485 ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2486 ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2487 ffi_1/nand_7/a Gnd 0.30fF
C2488 ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2489 ffi_1/qbar Gnd 0.60fF
C2490 ffi_1/nand_6/a Gnd 0.30fF
C2491 ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2492 ffi_1/inv_1/op Gnd 0.89fF
C2493 ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2494 ffi_1/nand_3/b Gnd 0.43fF
C2495 ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2496 ffi_1/nand_3/a Gnd 0.30fF
C2497 ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2498 ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2499 ffi_1/inv_0/op Gnd 0.26fF
C2500 ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2501 ffi_1/nand_1/a Gnd 0.30fF
C2502 ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2503 ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2504 ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2505 ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C2506 ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2507 ffipg_2/ffi_1/qbar Gnd 0.42fF
C2508 ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C2509 ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2510 ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C2511 ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2512 ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C2513 ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2514 ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C2515 ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2516 x3in Gnd 1.03fF
C2517 ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2518 ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C2519 ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2520 ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C2521 ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2522 ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2523 ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2524 ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C2525 ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2526 ffipg_2/ffi_0/qbar Gnd 0.42fF
C2527 ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C2528 ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2529 ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C2530 ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2531 ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C2532 ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2533 ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C2534 ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2535 y3in Gnd 1.03fF
C2536 ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2537 ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C2538 ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2539 ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C2540 ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2541 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2542 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2543 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2544 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2545 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2546 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2547 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2548 ffipg_2/ffi_0/q Gnd 2.68fF
C2549 ffipg_2/ffi_1/q Gnd 2.93fF
C2550 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2551 ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2552 ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2553 ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C2554 ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2555 ffipg_1/ffi_1/qbar Gnd 0.42fF
C2556 ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C2557 ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2558 ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C2559 ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2560 ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C2561 ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2562 ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C2563 ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2564 x2in Gnd 1.03fF
C2565 ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2566 ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C2567 ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2568 ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C2569 ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2570 ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2571 ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2572 ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C2573 ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2574 ffipg_1/ffi_0/qbar Gnd 0.42fF
C2575 ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C2576 ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2577 ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C2578 ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2579 ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C2580 ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2581 ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C2582 ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2583 y2in Gnd 0.94fF
C2584 ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2585 ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C2586 ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2587 ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C2588 ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2589 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2590 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2591 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2592 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2593 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2594 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2595 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2596 ffipg_1/ffi_0/q Gnd 2.68fF
C2597 ffipg_1/ffi_1/q Gnd 2.93fF
C2598 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2599 inv_9/in Gnd 0.23fF
C2600 nor_4/w_0_0# Gnd 1.81fF
C2601 ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2602 ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2603 ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C2604 ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2605 ffipg_0/ffi_1/qbar Gnd 0.42fF
C2606 ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C2607 ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2608 ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C2609 ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2610 ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C2611 ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2612 ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C2613 ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2614 x1in Gnd 0.91fF
C2615 ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2616 ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C2617 ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2618 ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C2619 ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2620 ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2621 ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2622 ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C2623 ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2624 ffipg_0/ffi_0/qbar Gnd 0.42fF
C2625 ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C2626 ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2627 ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C2628 ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2629 ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C2630 ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2631 ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C2632 ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2633 y1in Gnd 1.03fF
C2634 ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2635 ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C2636 ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2637 ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C2638 ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2639 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2640 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2641 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2642 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2643 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2644 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2645 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2646 ffipg_0/ffi_0/q Gnd 2.68fF
C2647 ffipg_0/ffi_1/q Gnd 2.93fF
C2648 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2649 nor_4/a Gnd 0.53fF
C2650 inv_8/in Gnd 0.22fF
C2651 inv_8/w_0_6# Gnd 1.40fF
C2652 inv_7/in Gnd 0.22fF
C2653 inv_7/w_0_6# Gnd 1.40fF
C2654 nor_4/b Gnd 0.22fF
C2655 nor_3/b Gnd 0.29fF
C2656 inv_5/in Gnd 0.22fF
C2657 inv_5/w_0_6# Gnd 1.40fF
C2658 cla_2/n Gnd 0.36fF
C2659 inv_6/in Gnd 0.23fF
C2660 nor_3/w_0_0# Gnd 1.81fF
C2661 cla_1/n Gnd 0.36fF
C2662 inv_4/in Gnd 0.23fF
C2663 nor_2/w_0_0# Gnd 1.81fF
C2664 cla_0/n Gnd 0.87fF
C2665 nor_2/b Gnd 0.88fF
C2666 inv_3/in Gnd 0.22fF
C2667 inv_3/w_0_6# Gnd 1.40fF
C2668 nor_1/b Gnd 0.68fF
C2669 inv_2/in Gnd 0.22fF
C2670 inv_2/w_0_6# Gnd 1.40fF
C2671 inv_1/in Gnd 0.23fF
C2672 nor_1/w_0_0# Gnd 1.81fF
C2673 inv_0/in Gnd 0.23fF
C2674 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C2675 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C2676 ffo_0/nand_7/a Gnd 0.30fF
C2677 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C2678 ffo_0/qbar Gnd 0.42fF
C2679 ffo_0/nand_6/a Gnd 0.30fF
C2680 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C2681 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C2682 ffo_0/nand_3/b Gnd 0.43fF
C2683 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C2684 ffo_0/nand_3/a Gnd 0.30fF
C2685 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C2686 ffo_0/nand_0/b Gnd 0.63fF
C2687 ffo_0/d Gnd 0.59fF
C2688 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C2689 ffo_0/inv_0/op Gnd 0.26fF
C2690 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C2691 ffo_0/nand_1/a Gnd 0.30fF
C2692 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C2693 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C2694 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C2695 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C2696 ffipg_3/k Gnd 2.02fF
C2697 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2698 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C2699 inv_4/op Gnd 1.37fF
C2700 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2701 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C2702 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C2703 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C2704 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C2705 sumffo_3/sbar Gnd 0.43fF
C2706 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C2707 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C2708 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C2709 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C2710 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C2711 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C2712 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C2713 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C2714 sumffo_3/ffo_0/d Gnd 0.64fF
C2715 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C2716 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C2717 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C2718 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C2719 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C2720 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C2721 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C2722 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C2723 nand_2/b Gnd 2.22fF
C2724 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2725 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C2726 ffipg_1/k Gnd 2.07fF
C2727 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2728 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C2729 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C2730 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C2731 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C2732 sumffo_1/sbar Gnd 0.43fF
C2733 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C2734 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C2735 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C2736 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C2737 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C2738 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C2739 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C2740 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C2741 sumffo_1/ffo_0/d Gnd 0.64fF
C2742 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C2743 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C2744 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C2745 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C2746 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C2747 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C2748 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C2749 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C2750 ffipg_2/k Gnd 2.04fF
C2751 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2752 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C2753 inv_1/op Gnd 1.37fF
C2754 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2755 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C2756 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C2757 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C2758 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C2759 sumffo_2/sbar Gnd 0.43fF
C2760 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C2761 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C2762 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C2763 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C2764 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C2765 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C2766 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C2767 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C2768 sumffo_2/ffo_0/d Gnd 0.64fF
C2769 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C2770 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C2771 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C2772 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C2773 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C2774 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C2775 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C2776 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C2777 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2778 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C2779 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2780 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C2781 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C2782 gnd Gnd 111.18fF
C2783 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C2784 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C2785 sumffo_0/sbar Gnd 0.43fF
C2786 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C2787 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C2788 clk Gnd 25.43fF
C2789 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C2790 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C2791 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C2792 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C2793 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C2794 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C2795 sumffo_0/ffo_0/d Gnd 0.64fF
C2796 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C2797 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C2798 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C2799 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C2800 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C2801 cla_2/p1 Gnd 1.09fF
C2802 cla_2/nor_1/w_0_0# Gnd 1.23fF
C2803 cla_2/nor_0/w_0_0# Gnd 1.23fF
C2804 cla_2/inv_0/in Gnd 0.27fF
C2805 cla_2/inv_0/w_0_6# Gnd 0.58fF
C2806 cla_2/g1 Gnd 0.45fF
C2807 cla_2/inv_0/op Gnd 0.26fF
C2808 cla_2/nand_0/w_0_0# Gnd 0.82fF
C2809 cla_1/nor_1/w_0_0# Gnd 1.23fF
C2810 cla_1/l Gnd 0.30fF
C2811 cla_1/nor_0/w_0_0# Gnd 1.23fF
C2812 cla_1/inv_0/in Gnd 0.27fF
C2813 cla_1/inv_0/w_0_6# Gnd 0.58fF
C2814 cla_1/inv_0/op Gnd 0.26fF
C2815 cla_1/nand_0/w_0_0# Gnd 0.82fF
C2816 inv_7/op Gnd 0.26fF
C2817 cla_0/nor_1/w_0_0# Gnd 1.23fF
C2818 cla_0/l Gnd 3.31fF
C2819 cla_0/nor_0/w_0_0# Gnd 1.23fF
C2820 cla_0/inv_0/in Gnd 0.27fF
C2821 cla_0/inv_0/w_0_6# Gnd 0.58fF
C2822 cla_0/inv_0/op Gnd 0.26fF
C2823 cla_0/nand_0/w_0_0# Gnd 0.82fF
C2824 cla_2/l Gnd 0.80fF
C2825 inv_0/op Gnd 0.23fF
C2826 nor_0/w_0_0# Gnd 2.63fF
C2827 ffipg_7/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2828 ffipg_7/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2829 ffipg_7/ffi_1/nand_7/a Gnd 0.30fF
C2830 ffipg_7/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2831 ffipg_7/ffi_1/qbar Gnd 0.42fF
C2832 ffipg_7/ffi_1/nand_6/a Gnd 0.30fF
C2833 ffipg_7/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2834 ffipg_7/ffi_1/inv_1/op Gnd 0.89fF
C2835 ffipg_7/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2836 ffipg_7/ffi_1/nand_3/b Gnd 0.43fF
C2837 ffipg_7/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2838 ffipg_7/ffi_1/nand_3/a Gnd 0.30fF
C2839 ffipg_7/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2840 ffipg_7/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2841 ffipg_7/ffi_1/inv_0/op Gnd 0.26fF
C2842 ffipg_7/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2843 ffipg_7/ffi_1/nand_1/a Gnd 0.30fF
C2844 ffipg_7/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2845 ffipg_7/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2846 ffipg_7/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2847 ffipg_7/ffi_0/nand_7/a Gnd 0.30fF
C2848 ffipg_7/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2849 ffipg_7/ffi_0/qbar Gnd 0.42fF
C2850 ffipg_7/ffi_0/nand_6/a Gnd 0.30fF
C2851 ffipg_7/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2852 ffipg_7/ffi_0/inv_1/op Gnd 0.89fF
C2853 ffipg_7/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2854 ffipg_7/ffi_0/nand_3/b Gnd 0.43fF
C2855 ffipg_7/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2856 ffipg_7/ffi_0/nand_3/a Gnd 0.30fF
C2857 ffipg_7/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2858 ffipg_7/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2859 ffipg_7/ffi_0/inv_0/op Gnd 0.26fF
C2860 ffipg_7/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2861 ffipg_7/ffi_0/nand_1/a Gnd 0.30fF
C2862 ffipg_7/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2863 ffipg_7/p Gnd 0.46fF
C2864 ffipg_7/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2865 ffipg_7/k Gnd 1.09fF
C2866 ffipg_7/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2867 ffipg_7/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2868 ffipg_7/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2869 ffipg_7/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2870 ffipg_7/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2871 ffipg_7/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2872 ffipg_7/g Gnd 0.16fF
C2873 ffipg_7/ffi_0/q Gnd 2.68fF
C2874 ffipg_7/ffi_1/q Gnd 2.93fF
C2875 ffipg_7/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2876 ffipg_6/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2877 ffipg_6/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2878 ffipg_6/ffi_1/nand_7/a Gnd 0.30fF
C2879 ffipg_6/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2880 ffipg_6/ffi_1/qbar Gnd 0.42fF
C2881 ffipg_6/ffi_1/nand_6/a Gnd 0.30fF
C2882 ffipg_6/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2883 ffipg_6/ffi_1/inv_1/op Gnd 0.89fF
C2884 ffipg_6/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2885 ffipg_6/ffi_1/nand_3/b Gnd 0.43fF
C2886 ffipg_6/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2887 ffipg_6/ffi_1/nand_3/a Gnd 0.30fF
C2888 ffipg_6/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2889 ffipg_6/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2890 ffipg_6/ffi_1/inv_0/op Gnd 0.26fF
C2891 ffipg_6/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2892 ffipg_6/ffi_1/nand_1/a Gnd 0.30fF
C2893 ffipg_6/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2894 ffipg_6/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2895 ffipg_6/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2896 ffipg_6/ffi_0/nand_7/a Gnd 0.30fF
C2897 ffipg_6/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2898 ffipg_6/ffi_0/qbar Gnd 0.42fF
C2899 ffipg_6/ffi_0/nand_6/a Gnd 0.30fF
C2900 ffipg_6/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2901 ffipg_6/ffi_0/inv_1/op Gnd 0.89fF
C2902 ffipg_6/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2903 ffipg_6/ffi_0/nand_3/b Gnd 0.43fF
C2904 ffipg_6/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2905 ffipg_6/ffi_0/nand_3/a Gnd 0.30fF
C2906 ffipg_6/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2907 ffipg_6/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2908 ffipg_6/ffi_0/inv_0/op Gnd 0.26fF
C2909 ffipg_6/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2910 ffipg_6/ffi_0/nand_1/a Gnd 0.30fF
C2911 ffipg_6/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2912 ffipg_6/p Gnd 0.46fF
C2913 ffipg_6/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2914 ffipg_6/k Gnd 1.09fF
C2915 ffipg_6/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2916 ffipg_6/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2917 ffipg_6/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2918 ffipg_6/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2919 ffipg_6/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2920 ffipg_6/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2921 ffipg_6/g Gnd 0.14fF
C2922 ffipg_6/ffi_0/q Gnd 2.68fF
C2923 ffipg_6/ffi_1/q Gnd 2.93fF
C2924 ffipg_6/pggen_0/nand_0/w_0_0# Gnd 0.82fF
