* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 vdd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 vdd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 s1 cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op s1 sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op s1 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 s1 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 vdd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 s3 ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op s3 sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op s3 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 s3 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 s2 nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op s2 sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op s2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 s2 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 vdd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 s4 ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op s4 sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op s4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 s4 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 vdd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in vdd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 vdd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in vdd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in vdd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 vdd y2in cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 cla_0/l x2in vdd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_0/l y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 vdd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in vdd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in vdd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 vdd y3in cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 cla_0/l x3in vdd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_0/l y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 vdd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in vdd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in vdd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 vdd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in vdd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 vdd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in vdd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in vdd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ffipg_1/pggen_0/xor_0/w_n3_4# gnd 0.02fF
C1 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C2 gnd cla_2/nand_0/a_13_n26# 0.01fF
C3 y4in cla_2/g1 0.13fF
C4 sumffo_3/xor_0/w_n3_4# inv_4/op 0.06fF
C5 gnd ffipg_0/k 0.41fF
C6 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C7 sumffo_1/xor_0/inv_0/w_0_6# vdd 0.09fF
C8 gnd y2in 1.68fF
C9 cla_2/l cla_0/n 0.32fF
C10 sumffo_1/xor_0/a_38_n43# cin 0.01fF
C11 ffipg_1/k cla_1/p0 0.05fF
C12 cla_2/p1 vdd 0.31fF
C13 cla_2/p0 cla_2/p1 0.24fF
C14 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.24fF
C15 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C16 cla_0/inv_0/w_0_6# vdd 0.06fF
C17 y4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C18 s2 sumffo_1/xor_0/a_10_10# 0.45fF
C19 gnd s2 0.14fF
C20 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C21 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/k 0.21fF
C22 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C23 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C24 nor_0/a gnd 0.23fF
C25 nor_2/w_0_0# inv_4/in 0.11fF
C26 gnd cla_2/l 0.24fF
C27 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C28 sumffo_3/xor_0/inv_1/op vdd 0.15fF
C29 sumffo_3/xor_0/w_n3_4# cin 0.01fF
C30 inv_2/in inv_2/w_0_6# 0.10fF
C31 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C32 gnd y1in 1.62fF
C33 nor_4/a nor_4/b 0.42fF
C34 gnd s1 0.14fF
C35 cla_0/g0 vdd 0.53fF
C36 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C37 ffipg_0/k sumffo_0/xor_0/w_n3_4# 0.06fF
C38 nor_0/w_0_0# cin 0.16fF
C39 inv_2/w_0_6# nand_2/b 0.03fF
C40 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C41 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C42 inv_9/in vdd 0.09fF
C43 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C44 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C45 cla_2/inv_0/in cla_2/p1 0.02fF
C46 y4in ffipg_3/k 0.07fF
C47 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C48 nor_2/b inv_3/in 0.04fF
C49 ffipg_3/k sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C50 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C51 nor_3/b cla_2/n 0.41fF
C52 inv_5/in cla_2/l 0.05fF
C53 ffipg_1/k gnd 0.39fF
C54 ffipg_0/pggen_0/nor_0/w_0_0# y1in 0.06fF
C55 ffipg_3/k x4in 0.46fF
C56 sumffo_2/xor_0/a_10_10# cin 0.04fF
C57 gnd inv_7/op 0.10fF
C58 inv_1/op gnd 0.32fF
C59 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C60 s4 cin 0.16fF
C61 s3 cin 0.28fF
C62 ffipg_2/pggen_0/xor_0/w_n3_4# y3in 0.06fF
C63 vdd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C64 sumffo_2/xor_0/a_10_10# ffipg_2/k 0.12fF
C65 cla_0/l cla_2/p1 0.30fF
C66 inv_0/op cla_0/g0 0.32fF
C67 y4in ffipg_3/pggen_0/xor_0/inv_0/op 0.20fF
C68 y1in ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C69 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C70 sumffo_0/xor_0/w_n3_4# s1 0.02fF
C71 cla_2/nor_0/w_0_0# vdd 0.31fF
C72 cla_1/inv_0/op vdd 0.17fF
C73 cla_0/inv_0/op nand_2/b 0.09fF
C74 vdd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C75 ffipg_1/pggen_0/nand_0/w_0_0# y2in 0.06fF
C76 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C77 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C78 ffipg_2/pggen_0/xor_0/inv_1/op x3in 0.06fF
C79 ffipg_3/pggen_0/xor_0/inv_0/op x4in 0.27fF
C80 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C81 ffipg_0/k cin 0.19fF
C82 ffipg_2/pggen_0/nor_0/w_0_0# x3in 0.06fF
C83 gnd x1in 0.22fF
C84 cla_0/l cla_0/g0 0.14fF
C85 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C86 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# x4in 0.06fF
C87 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C88 x1in ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C89 cla_0/nor_1/w_0_0# vdd 0.31fF
C90 inv_5/w_0_6# vdd 0.15fF
C91 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.21fF
C92 cin sumffo_0/xor_0/a_10_10# 0.12fF
C93 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k 0.06fF
C94 s2 cin 0.27fF
C95 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C96 sumffo_3/xor_0/a_10_10# cin 0.04fF
C97 nor_3/w_0_0# vdd 0.14fF
C98 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k 0.52fF
C99 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C100 cla_1/n vdd 0.28fF
C101 cla_1/p0 cla_0/g0 0.38fF
C102 ffipg_0/pggen_0/nor_0/w_0_0# x1in 0.06fF
C103 cla_2/p0 vdd 0.43fF
C104 inv_0/in vdd 0.07fF
C105 nor_3/w_0_0# inv_6/in 0.11fF
C106 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C107 inv_6/in vdd 0.09fF
C108 gnd cla_2/p1 0.68fF
C109 s3 sumffo_2/xor_0/inv_1/op 0.52fF
C110 x2in ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C111 ffipg_0/pggen_0/xor_0/inv_0/op y1in 0.20fF
C112 cla_1/inv_0/op cla_0/l 0.35fF
C113 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C114 ffipg_1/k cin 0.06fF
C115 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C116 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C117 inv_7/op cin 0.31fF
C118 inv_0/op vdd 0.17fF
C119 sumffo_3/xor_0/inv_1/op gnd 0.20fF
C120 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C121 inv_0/op inv_0/in 0.04fF
C122 inv_7/op inv_8/w_0_6# 0.06fF
C123 cla_2/inv_0/in vdd 0.05fF
C124 inv_1/op ffipg_2/k 0.09fF
C125 gnd cla_0/g0 0.70fF
C126 cla_1/l vdd 0.22fF
C127 inv_9/in cout 0.04fF
C128 cla_2/p0 cla_1/l 0.02fF
C129 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C130 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C131 sumffo_1/xor_0/inv_0/op cin 0.06fF
C132 gnd inv_9/in 0.24fF
C133 nor_1/b vdd 0.25fF
C134 sumffo_0/xor_0/inv_1/op vdd 0.15fF
C135 cla_0/l cla_1/n 0.13fF
C136 cla_0/nand_0/w_0_0# vdd 0.10fF
C137 cla_0/l vdd 1.60fF
C138 cla_2/p0 cla_0/l 0.44fF
C139 inv_3/w_0_6# vdd 0.15fF
C140 cla_1/inv_0/op cla_0/n 0.06fF
C141 ffipg_3/pggen_0/xor_0/inv_1/op vdd 0.15fF
C142 cla_1/p0 cla_0/nor_1/w_0_0# 0.06fF
C143 vdd ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C144 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C145 nor_3/b cla_2/l 0.10fF
C146 sumffo_2/xor_0/w_n3_4# s3 0.02fF
C147 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C148 cla_1/p0 vdd 0.43fF
C149 cla_2/p0 cla_1/p0 0.24fF
C150 ffipg_3/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C151 inv_1/op nor_1/w_0_0# 0.03fF
C152 sumffo_1/xor_0/w_n3_4# s2 0.02fF
C153 gnd cla_1/inv_0/op 0.10fF
C154 x1in ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C155 inv_7/w_0_6# inv_7/in 0.10fF
C156 nor_0/w_0_0# nand_2/b 0.04fF
C157 inv_5/w_0_6# cla_0/n 0.06fF
C158 sumffo_3/xor_0/inv_1/op inv_4/op 0.06fF
C159 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C160 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C161 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C162 cla_2/inv_0/in cla_0/l 0.16fF
C163 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C164 cla_2/nor_1/w_0_0# vdd 0.31fF
C165 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C166 cla_0/n vdd 0.56fF
C167 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C168 inv_9/in nor_4/a 0.02fF
C169 cla_0/l cla_1/l 0.08fF
C170 y4in ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C171 cla_1/l inv_3/w_0_6# 0.06fF
C172 gnd inv_5/w_0_6# 0.26fF
C173 sumffo_1/xor_0/inv_1/op s2 0.52fF
C174 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C175 cla_1/nand_0/w_0_0# vdd 0.10fF
C176 cla_2/g1 cla_2/n 0.13fF
C177 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C178 cla_0/nand_0/w_0_0# cla_0/l 0.06fF
C179 vdd cout 0.15fF
C180 sumffo_3/xor_0/inv_1/op cin 0.04fF
C181 gnd cla_1/n 0.24fF
C182 sumffo_1/xor_0/a_10_10# vdd 0.93fF
C183 gnd vdd 3.73fF
C184 gnd cla_2/p0 0.68fF
C185 cla_1/p0 cla_1/l 0.16fF
C186 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# x3in 0.06fF
C187 gnd inv_0/in 0.24fF
C188 y1in ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C189 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C190 vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C191 cla_0/g0 cin 0.08fF
C192 gnd inv_6/in 0.24fF
C193 inv_5/in inv_5/w_0_6# 0.10fF
C194 cla_0/l cla_1/p0 0.09fF
C195 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C196 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C197 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C198 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C199 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_0/op 0.06fF
C200 inv_8/in vdd 0.30fF
C201 ffipg_0/pggen_0/nor_0/w_0_0# vdd 0.11fF
C202 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C203 cla_1/l cla_0/n 0.07fF
C204 inv_5/in vdd 0.30fF
C205 nor_2/b nor_2/w_0_0# 0.06fF
C206 x3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C207 sumffo_2/xor_0/inv_0/op s3 0.06fF
C208 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C209 inv_1/op inv_1/in 0.04fF
C210 gnd inv_0/op 0.10fF
C211 sumffo_2/xor_0/w_n3_4# inv_1/op 0.06fF
C212 nor_1/b cla_0/n 0.36fF
C213 ffipg_2/pggen_0/xor_0/inv_0/op vdd 0.15fF
C214 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C215 cla_2/inv_0/in gnd 0.30fF
C216 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C217 cla_0/l cla_0/n 0.25fF
C218 sumffo_0/xor_0/w_n3_4# vdd 0.12fF
C219 inv_3/w_0_6# cla_0/n 0.16fF
C220 y4in cla_2/p1 0.03fF
C221 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C222 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_0/op 0.08fF
C223 sumffo_2/xor_0/inv_0/w_0_6# vdd 0.09fF
C224 gnd cla_1/l 0.18fF
C225 vdd ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C226 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_1/w_0_6# 0.03fF
C227 cla_1/nand_0/w_0_0# cla_0/l 0.06fF
C228 x4in cla_2/p1 0.22fF
C229 ffipg_1/pggen_0/xor_0/w_n3_4# x2in 0.06fF
C230 nor_4/a vdd 0.19fF
C231 cla_2/inv_0/op vdd 0.17fF
C232 gnd nor_1/b 0.10fF
C233 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C234 y4in ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C235 gnd cla_0/nand_0/w_0_0# 0.01fF
C236 inv_7/in inv_7/op 0.04fF
C237 inv_4/op vdd 0.26fF
C238 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C239 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_1/w_0_6# 0.03fF
C240 ffipg_1/k nand_2/b 0.15fF
C241 gnd cla_0/l 1.69fF
C242 gnd inv_3/w_0_6# 0.02fF
C243 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C244 ffipg_0/pggen_0/nand_0/a_13_n26# vdd 0.01fF
C245 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.24fF
C246 y2in x2in 0.73fF
C247 x3in vdd 0.93fF
C248 cla_2/p0 x3in 0.22fF
C249 cla_1/inv_0/w_0_6# vdd 0.06fF
C250 ffipg_1/pggen_0/nand_0/w_0_0# vdd 0.10fF
C251 gnd cla_1/p0 0.68fF
C252 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C253 ffipg_3/k sumffo_3/xor_0/inv_0/op 0.20fF
C254 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C255 sumffo_1/xor_0/inv_1/w_0_6# nand_2/b 0.23fF
C256 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/k 0.01fF
C257 cin vdd 0.78fF
C258 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C259 vdd ffipg_1/pggen_0/nand_0/a_13_n26# 0.01fF
C260 inv_0/in cin 0.07fF
C261 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C262 inv_8/w_0_6# vdd 0.15fF
C263 ffipg_2/k vdd 0.35fF
C264 cla_2/p0 ffipg_2/k 0.05fF
C265 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C266 gnd cla_0/n 0.61fF
C267 ffipg_2/pggen_0/xor_0/a_10_10# vdd 0.93fF
C268 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C269 ffipg_0/pggen_0/xor_0/inv_0/op vdd 0.15fF
C270 gnd cla_1/nand_0/w_0_0# 0.01fF
C271 ffipg_1/k x2in 0.46fF
C272 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C273 cla_2/nand_0/w_0_0# vdd 0.10fF
C274 cla_1/n inv_4/in 0.02fF
C275 gnd cout 0.10fF
C276 vdd inv_4/in 0.09fF
C277 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C278 ffipg_2/pggen_0/nand_0/a_13_n26# vdd 0.01fF
C279 inv_5/in cla_0/n 0.13fF
C280 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C281 nor_0/a cla_0/nor_0/w_0_0# 0.06fF
C282 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C283 ffipg_2/pggen_0/xor_0/inv_1/op y3in 0.22fF
C284 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C285 sumffo_0/xor_0/inv_0/op s1 0.06fF
C286 gnd inv_8/in 0.13fF
C287 nor_1/w_0_0# vdd 0.17fF
C288 ffipg_1/pggen_0/xor_0/a_10_10# y2in 0.12fF
C289 ffipg_2/pggen_0/nor_0/w_0_0# y3in 0.06fF
C290 sumffo_0/xor_0/inv_1/op cin 0.22fF
C291 nor_3/b inv_5/w_0_6# 0.17fF
C292 gnd inv_5/in 0.19fF
C293 cla_0/l cin 0.33fF
C294 y4in vdd 0.10fF
C295 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C296 sumffo_3/xor_0/inv_1/w_0_6# vdd 0.06fF
C297 x4in vdd 0.93fF
C298 nor_3/b nor_3/w_0_0# 0.06fF
C299 s4 sumffo_3/xor_0/inv_0/op 0.06fF
C300 cla_0/l ffipg_2/k 0.10fF
C301 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.21fF
C302 sumffo_2/xor_0/inv_1/op vdd 0.15fF
C303 nor_3/b vdd 0.23fF
C304 x2in ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C305 s4 sumffo_3/xor_0/w_n3_4# 0.02fF
C306 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C307 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C308 cla_0/g0 nand_2/b 0.13fF
C309 nor_4/b nor_4/w_0_0# 0.06fF
C310 cla_1/p0 ffipg_2/k 0.06fF
C311 gnd nor_4/a 0.21fF
C312 nor_3/b inv_6/in 0.16fF
C313 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C314 gnd cla_2/inv_0/op 0.10fF
C315 cinbar nor_0/w_0_0# 0.06fF
C316 gnd inv_4/op 0.32fF
C317 sumffo_1/xor_0/w_n3_4# vdd 0.12fF
C318 inv_3/in vdd 0.30fF
C319 gnd x3in 0.31fF
C320 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/k 0.45fF
C321 cla_1/nor_1/w_0_0# vdd 0.31fF
C322 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C323 nor_4/a inv_8/in 0.04fF
C324 sumffo_2/xor_0/a_10_10# s3 0.45fF
C325 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C326 nor_1/w_0_0# nor_1/b 0.06fF
C327 ffipg_2/k cla_0/n 0.06fF
C328 ffipg_2/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C329 sumffo_1/xor_0/inv_1/op vdd 0.15fF
C330 sumffo_1/xor_0/a_10_10# cin 0.06fF
C331 gnd cin 0.74fF
C332 y4in ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C333 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C334 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C335 inv_1/in vdd 0.09fF
C336 sumffo_2/xor_0/w_n3_4# vdd 0.12fF
C337 vdd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C338 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C339 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C340 gnd ffipg_2/k 0.29fF
C341 cinbar ffipg_0/k 0.06fF
C342 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C343 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C344 ffipg_2/pggen_0/xor_0/inv_0/op x3in 0.27fF
C345 inv_2/in vdd 0.30fF
C346 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.17fF
C347 y4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C348 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C349 inv_8/in cin 0.13fF
C350 cla_2/g1 cla_2/p1 0.00fF
C351 cla_2/nand_0/w_0_0# gnd 0.08fF
C352 x4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C353 nor_0/a nor_0/w_0_0# 0.06fF
C354 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C355 inv_8/in inv_8/w_0_6# 0.10fF
C356 gnd inv_4/in 0.24fF
C357 inv_7/in vdd 0.30fF
C358 cla_0/g0 cla_0/inv_0/in 0.16fF
C359 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C360 inv_7/w_0_6# cla_2/l 0.06fF
C361 nor_1/w_0_0# cla_0/n 0.06fF
C362 nor_0/a cinbar 0.32fF
C363 nand_2/b vdd 0.92fF
C364 x2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C365 inv_3/w_0_6# inv_3/in 0.10fF
C366 sumffo_3/xor_0/a_10_10# s4 0.45fF
C367 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C368 sumffo_0/xor_0/w_n3_4# cin 0.06fF
C369 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C370 ffipg_1/pggen_0/xor_0/w_n3_4# y2in 0.06fF
C371 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C372 sumffo_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C373 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C374 cla_1/inv_0/in vdd 0.05fF
C375 cla_2/p0 cla_1/inv_0/in 0.02fF
C376 inv_1/in nor_1/b 0.16fF
C377 nor_4/a inv_8/w_0_6# 0.03fF
C378 y4in gnd 1.66fF
C379 inv_7/w_0_6# inv_7/op 0.03fF
C380 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C381 gnd x4in 0.31fF
C382 cla_2/inv_0/w_0_6# vdd 0.06fF
C383 gnd cla_1/nand_0/a_13_n26# 0.01fF
C384 nor_0/a ffipg_0/k 0.05fF
C385 y1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C386 inv_2/in nor_1/b 0.04fF
C387 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C388 gnd nor_3/b 0.10fF
C389 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# y1in 0.23fF
C390 ffipg_2/k x3in 0.46fF
C391 ffipg_0/k y1in 0.07fF
C392 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C393 ffipg_3/k cla_2/p1 0.05fF
C394 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C395 sumffo_2/xor_0/inv_0/op vdd 0.15fF
C396 nand_2/b cla_1/l 0.31fF
C397 inv_2/w_0_6# vdd 0.15fF
C398 x2in vdd 0.93fF
C399 inv_4/op inv_4/in 0.04fF
C400 y1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C401 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/k 0.02fF
C402 cla_0/l inv_7/in 0.13fF
C403 sumffo_0/xor_0/inv_1/w_0_6# vdd 0.07fF
C404 sumffo_3/xor_0/inv_1/op ffipg_3/k 0.22fF
C405 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C406 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C407 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C408 cla_0/l nand_2/b 0.06fF
C409 inv_8/w_0_6# cin 0.06fF
C410 s1 sumffo_0/xor_0/a_10_10# 0.45fF
C411 nand_2/b inv_3/w_0_6# 0.06fF
C412 gnd inv_3/in 0.17fF
C413 nor_0/a y1in 0.03fF
C414 gnd cla_0/nand_0/a_13_n26# 0.00fF
C415 nor_3/b inv_5/in 0.04fF
C416 ffipg_1/k y2in 0.07fF
C417 inv_1/in cla_0/n 0.02fF
C418 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C419 sumffo_2/xor_0/inv_1/w_0_6# vdd 0.06fF
C420 cla_0/inv_0/in vdd 0.05fF
C421 ffipg_3/pggen_0/nand_0/w_0_0# vdd 0.10fF
C422 y3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C423 cla_0/l cla_1/inv_0/in 0.23fF
C424 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C425 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C426 cla_0/inv_0/op vdd 0.17fF
C427 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C428 ffipg_1/k nor_0/a 0.06fF
C429 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C430 vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C431 gnd inv_1/in 0.24fF
C432 cla_2/g1 vdd 0.35fF
C433 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C434 sumffo_0/xor_0/inv_0/op vdd 0.15fF
C435 x1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C436 cla_0/nor_0/w_0_0# vdd 0.31fF
C437 nand_2/b cla_0/n 0.06fF
C438 inv_2/w_0_6# nor_1/b 0.03fF
C439 sumffo_1/xor_0/inv_0/op s2 0.06fF
C440 gnd inv_2/in 0.17fF
C441 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C442 x1in ffipg_0/k 0.46fF
C443 inv_2/w_0_6# cla_0/l 0.06fF
C444 vdd y3in 0.15fF
C445 nor_2/b cla_1/n 0.39fF
C446 cla_2/p0 y3in 0.03fF
C447 inv_9/in nor_4/w_0_0# 0.11fF
C448 nor_2/b vdd 0.21fF
C449 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C450 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C451 ffipg_3/pggen_0/nor_0/w_0_0# vdd 0.11fF
C452 x2in ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C453 gnd inv_7/in 0.13fF
C454 x1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C455 y2in ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C456 sumffo_3/xor_0/inv_0/w_0_6# vdd 0.09fF
C457 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C458 gnd nand_2/b 0.94fF
C459 cin sumffo_2/xor_0/inv_1/op 0.04fF
C460 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C461 cla_0/g0 nor_0/w_0_0# 0.06fF
C462 cla_1/p0 x2in 0.22fF
C463 nor_0/a x1in 0.22fF
C464 nor_3/w_0_0# cla_2/n 0.06fF
C465 cla_2/inv_0/in cla_2/g1 0.04fF
C466 ffipg_1/pggen_0/xor_0/a_10_10# vdd 0.93fF
C467 sumffo_3/xor_0/inv_1/op s4 0.52fF
C468 cla_0/l cla_0/inv_0/in 0.07fF
C469 gnd sumffo_0/xor_0/inv_0/w_0_6# 0.02fF
C470 sumffo_2/xor_0/a_38_n43# cin 0.01fF
C471 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C472 x1in y1in 0.73fF
C473 vdd cla_2/n 0.28fF
C474 gnd cla_1/inv_0/in 0.30fF
C475 ffipg_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C476 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C477 cla_0/l cla_0/inv_0/op 0.35fF
C478 ffipg_2/pggen_0/xor_0/w_n3_4# x3in 0.06fF
C479 sumffo_1/xor_0/w_n3_4# cin 0.00fF
C480 ffipg_3/k vdd 0.35fF
C481 ffipg_3/k cla_2/p0 0.06fF
C482 inv_6/in cla_2/n 0.02fF
C483 cla_1/p0 cla_0/inv_0/in 0.02fF
C484 cla_0/l cla_2/g1 0.26fF
C485 cla_1/n nor_2/w_0_0# 0.06fF
C486 nor_2/w_0_0# vdd 0.17fF
C487 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C488 inv_9/in nor_4/b 0.16fF
C489 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C490 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C491 cla_2/l cla_2/p1 0.02fF
C492 gnd inv_2/w_0_6# 0.02fF
C493 sumffo_2/xor_0/inv_0/op gnd 0.17fF
C494 cla_0/l y3in 0.13fF
C495 sumffo_1/xor_0/inv_1/op cin 0.04fF
C496 gnd x2in 0.31fF
C497 nor_2/b inv_3/w_0_6# 0.03fF
C498 ffipg_3/pggen_0/xor_0/inv_0/op vdd 0.15fF
C499 sumffo_3/xor_0/inv_0/op vdd 0.15fF
C500 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C501 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C502 sumffo_2/xor_0/w_n3_4# cin 0.00fF
C503 y4in x4in 0.73fF
C504 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C505 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C506 vdd nor_4/w_0_0# 0.15fF
C507 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C508 sumffo_3/xor_0/w_n3_4# vdd 0.12fF
C509 ffipg_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C510 sumffo_2/xor_0/w_n3_4# ffipg_2/k 0.06fF
C511 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C512 inv_2/in cin 0.13fF
C513 nor_0/a cla_0/g0 0.57fF
C514 gnd cla_0/inv_0/in 0.30fF
C515 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C516 cla_0/g0 y1in 0.13fF
C517 gnd cla_0/inv_0/op 0.10fF
C518 y2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C519 nor_0/w_0_0# vdd 0.46fF
C520 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C521 nor_0/w_0_0# inv_0/in 0.11fF
C522 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C523 ffipg_3/k cla_0/l 0.10fF
C524 inv_7/w_0_6# vdd 0.15fF
C525 nand_2/b cin 0.04fF
C526 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C527 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C528 cinbar vdd 0.16fF
C529 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C530 gnd cla_2/g1 0.30fF
C531 sumffo_2/xor_0/a_10_10# vdd 0.93fF
C532 cinbar inv_0/in 0.16fF
C533 gnd sumffo_0/xor_0/inv_0/op 0.21fF
C534 ffipg_2/k nand_2/b 0.06fF
C535 nor_3/w_0_0# nor_4/b 0.03fF
C536 ffipg_1/k cla_0/g0 0.06fF
C537 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C538 nor_4/b vdd 0.15fF
C539 nor_1/w_0_0# inv_1/in 0.11fF
C540 gnd y3in 1.68fF
C541 gnd nor_2/b 0.10fF
C542 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C543 inv_0/op nor_0/w_0_0# 0.10fF
C544 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C545 ffipg_1/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C546 ffipg_0/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C547 nor_4/b inv_6/in 0.04fF
C548 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C549 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C550 ffipg_1/pggen_0/nand_0/w_0_0# x2in 0.06fF
C551 ffipg_0/k vdd 0.33fF
C552 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C553 ffipg_3/k cla_0/n 0.06fF
C554 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C555 y2in vdd 0.15fF
C556 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C557 sumffo_3/xor_0/a_38_n43# cin 0.01fF
C558 sumffo_2/xor_0/inv_0/op cin 0.06fF
C559 inv_2/w_0_6# cin 0.06fF
C560 gnd cla_2/n 0.32fF
C561 vdd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C562 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C563 inv_5/w_0_6# cla_2/l 0.08fF
C564 ffipg_2/pggen_0/xor_0/inv_1/op vdd 0.15fF
C565 sumffo_0/xor_0/a_10_10# vdd 0.93fF
C566 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C567 sumffo_3/xor_0/a_10_10# vdd 0.93fF
C568 cla_1/nor_0/w_0_0# vdd 0.31fF
C569 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C570 sumffo_0/xor_0/inv_1/w_0_6# cin 0.23fF
C571 cla_2/g1 cla_2/inv_0/op 0.35fF
C572 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C573 inv_7/w_0_6# cla_0/l 0.06fF
C574 ffipg_3/k gnd 0.31fF
C575 ffipg_2/pggen_0/xor_0/inv_0/op y3in 0.20fF
C576 nor_0/a vdd 0.35fF
C577 ffipg_2/pggen_0/nor_0/w_0_0# vdd 0.11fF
C578 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C579 cla_2/p0 cla_2/l 0.16fF
C580 cla_2/l vdd 0.38fF
C581 nor_0/a inv_0/in 0.02fF
C582 y1in vdd 0.15fF
C583 sumffo_2/xor_0/inv_1/w_0_6# ffipg_2/k 0.23fF
C584 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.21fF
C585 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C586 ffipg_1/k vdd 0.36fF
C587 x3in y3in 0.73fF
C588 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C589 nor_4/w_0_0# cout 0.03fF
C590 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C591 inv_1/op vdd 0.26fF
C592 inv_7/op vdd 0.17fF
C593 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C594 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C595 sumffo_0/xor_0/inv_0/op cin 0.20fF
C596 nand_2/b inv_3/in 0.13fF
C597 cla_0/l y2in 0.13fF
C598 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C599 y2in ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C600 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.02fF
C601 ffipg_3/pggen_0/xor_0/a_10_10# vdd 0.93fF
C602 sumffo_1/xor_0/inv_0/op vdd 0.15fF
C603 sumffo_1/xor_0/inv_1/w_0_6# vdd 0.06fF
C604 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C605 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C606 ffipg_3/k inv_4/op 0.09fF
C607 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C608 cla_1/p0 y2in 0.03fF
C609 sumffo_1/xor_0/inv_1/op nand_2/b 0.22fF
C610 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C611 nor_0/a cla_0/l 0.16fF
C612 ffipg_2/k y3in 0.07fF
C613 cla_0/l cla_2/l 0.37fF
C614 inv_4/op nor_2/w_0_0# 0.03fF
C615 ffipg_2/pggen_0/xor_0/a_10_10# y3in 0.12fF
C616 sumffo_0/xor_0/inv_1/op s1 0.52fF
C617 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C618 x1in vdd 0.97fF
C619 gnd s4 0.14fF
C620 gnd s3 0.14fF
C621 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C622 y4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C623 nor_0/a cla_1/p0 0.24fF
C624 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C625 inv_2/in nand_2/b 0.34fF
C626 gnd nor_4/b 0.10fF
C627 vdd ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C628 nor_2/b inv_4/in 0.16fF
C629 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C630 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C631 y2in ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C632 nor_4/a nor_4/w_0_0# 0.07fF
C633 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C634 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C635 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C636 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C637 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C638 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C639 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C640 y4in Gnd 2.72fF
C641 x4in Gnd 2.80fF
C642 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C643 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C644 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C645 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C646 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C647 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C648 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C649 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C650 y3in Gnd 2.72fF
C651 x3in Gnd 2.80fF
C652 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C653 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C654 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C655 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C656 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C657 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C658 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C659 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C660 y2in Gnd 2.72fF
C661 x2in Gnd 2.80fF
C662 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C663 cout Gnd 0.19fF
C664 inv_9/in Gnd 0.23fF
C665 nor_4/w_0_0# Gnd 1.81fF
C666 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C667 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C668 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C669 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C670 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C671 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C672 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C673 y1in Gnd 2.72fF
C674 x1in Gnd 2.80fF
C675 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C676 nor_4/a Gnd 0.59fF
C677 inv_8/in Gnd 0.22fF
C678 inv_8/w_0_6# Gnd 1.40fF
C679 inv_7/in Gnd 0.22fF
C680 inv_7/w_0_6# Gnd 1.40fF
C681 nor_4/b Gnd 0.32fF
C682 nor_3/b Gnd 0.77fF
C683 inv_5/in Gnd 0.22fF
C684 inv_5/w_0_6# Gnd 1.40fF
C685 cla_2/n Gnd 0.36fF
C686 inv_6/in Gnd 0.23fF
C687 nor_3/w_0_0# Gnd 1.81fF
C688 vdd Gnd 8.88fF
C689 cla_1/n Gnd 0.36fF
C690 inv_4/in Gnd 0.23fF
C691 nor_2/w_0_0# Gnd 1.81fF
C692 cla_0/n Gnd 1.34fF
C693 nor_2/b Gnd 0.82fF
C694 inv_3/in Gnd 0.22fF
C695 inv_3/w_0_6# Gnd 1.40fF
C696 cinbar Gnd 1.21fF
C697 nor_0/a Gnd 2.07fF
C698 nor_1/b Gnd 1.05fF
C699 inv_2/in Gnd 0.22fF
C700 inv_2/w_0_6# Gnd 1.40fF
C701 inv_1/in Gnd 0.23fF
C702 nor_1/w_0_0# Gnd 1.81fF
C703 inv_0/in Gnd 0.23fF
C704 s4 Gnd 0.07fF
C705 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C706 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C707 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C708 ffipg_3/k Gnd 2.89fF
C709 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C710 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C711 inv_4/op Gnd 1.37fF
C712 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C713 s2 Gnd 0.07fF
C714 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C715 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C716 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C717 nand_2/b Gnd 2.36fF
C718 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C719 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C720 ffipg_1/k Gnd 2.78fF
C721 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C722 s3 Gnd 0.07fF
C723 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C724 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C725 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C726 ffipg_2/k Gnd 2.89fF
C727 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C728 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C729 inv_1/op Gnd 1.30fF
C730 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C731 s1 Gnd 0.07fF
C732 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C733 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C734 gnd Gnd 23.13fF
C735 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C736 cin Gnd 7.80fF
C737 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C738 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C739 ffipg_0/k Gnd 1.49fF
C740 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C741 cla_2/p1 Gnd 1.09fF
C742 cla_2/nor_1/w_0_0# Gnd 1.23fF
C743 cla_2/nor_0/w_0_0# Gnd 1.23fF
C744 cla_2/inv_0/in Gnd 0.27fF
C745 cla_2/inv_0/w_0_6# Gnd 0.58fF
C746 cla_2/g1 Gnd 0.59fF
C747 cla_2/inv_0/op Gnd 0.26fF
C748 cla_2/nand_0/w_0_0# Gnd 0.82fF
C749 cla_2/p0 Gnd 0.38fF
C750 cla_1/nor_1/w_0_0# Gnd 1.23fF
C751 cla_1/l Gnd 0.30fF
C752 cla_1/nor_0/w_0_0# Gnd 1.23fF
C753 cla_1/inv_0/in Gnd 0.27fF
C754 cla_1/inv_0/w_0_6# Gnd 0.58fF
C755 cla_1/inv_0/op Gnd 0.26fF
C756 cla_1/nand_0/w_0_0# Gnd 0.82fF
C757 inv_7/op Gnd 0.26fF
C758 cla_1/p0 Gnd 2.28fF
C759 cla_0/nor_1/w_0_0# Gnd 1.23fF
C760 cla_0/l Gnd 3.41fF
C761 cla_0/nor_0/w_0_0# Gnd 1.23fF
C762 cla_0/inv_0/in Gnd 0.27fF
C763 cla_0/inv_0/w_0_6# Gnd 0.58fF
C764 cla_0/inv_0/op Gnd 0.26fF
C765 cla_0/nand_0/w_0_0# Gnd 0.82fF
C766 cla_2/l Gnd 0.25fF
C767 cla_0/g0 Gnd 1.40fF
C768 inv_0/op Gnd 0.23fF
C769 nor_0/w_0_0# Gnd 2.63fF
