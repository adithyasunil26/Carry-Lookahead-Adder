* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0

M1004 vdd b a_10_10# w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1005 op b a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1006 gnd inv_1/op a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1007 a_10_10# inv_1/op op w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1008 a_10_n43# a gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_38_n43# inv_0/op op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_10_10# a vdd w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 op inv_0/op a_10_10# w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 inv_0/op inv_1/op 0.08fF
C1 a b 0.09fF
C2 a_10_10# b 0.12fF
C3 w_n3_4# b 0.06fF
C4 gnd b 0.11fF
C5 a inv_1/op 0.06fF
C6 w_n3_4# inv_1/op 0.06fF
C7 inv_0/op a 0.27fF
C8 w_n3_4# inv_0/op 0.06fF
C9 inv_1/op gnd 0.20fF
C10 inv_0/op inv_0/w_0_6# 0.03fF
C11 vdd b 0.10fF
C12 inv_0/op gnd 0.17fF
C13 w_n3_4# a 0.06fF
C14 vdd inv_1/w_0_6# 0.06fF
C15 inv_1/op op 0.52fF
C16 w_n3_4# a_10_10# 0.16fF
C17 inv_1/op vdd 0.15fF
C18 a inv_0/w_0_6# 0.06fF
C19 inv_0/op op 0.06fF
C20 inv_0/op vdd 0.15fF
C21 a gnd 0.22fF
C22 inv_1/w_0_6# b 0.23fF
C23 inv_1/op b 0.22fF
C24 a vdd 0.11fF
C25 a_10_10# op 0.45fF
C26 w_n3_4# op 0.02fF
C27 vdd a_10_10# 0.93fF
C28 w_n3_4# vdd 0.12fF
C29 inv_0/op b 0.20fF
C30 inv_0/w_0_6# vdd 0.09fF
C31 inv_1/op inv_1/w_0_6# 0.03fF
C32 gnd op 0.14fF
C33 gnd vdd 0.25fF
C34 op Gnd 0.04fF
C35 a_10_10# Gnd 0.01fF
C36 w_n3_4# Gnd 1.14fF
C37 gnd Gnd 0.72fF
C38 inv_1/op Gnd 0.49fF
C39 vdd Gnd 0.59fF
C40 b Gnd 1.37fF
C41 inv_1/w_0_6# Gnd 0.58fF
C42 inv_0/op Gnd 0.50fF
C43 a Gnd 1.28fF
C44 inv_0/w_0_6# Gnd 0.58fF
