magic
tech scmos
timestamp 1619200732
<< metal1 >>
rect -3 1270 97 1273
rect 102 1270 546 1273
rect 3 1263 410 1266
rect 3 1256 6 1263
rect -3 1252 0 1255
rect 241 1212 260 1215
rect 233 1183 244 1186
rect 241 1156 254 1159
rect -3 1153 0 1156
rect -3 1083 0 1086
rect 251 1047 254 1156
rect 257 1056 260 1212
rect 278 1145 293 1148
rect 278 1054 281 1145
rect 415 1143 418 1146
rect 641 1137 644 1140
rect 262 1051 281 1054
rect 251 1044 497 1047
rect 479 1014 484 1019
rect 494 998 497 1044
rect 539 1026 542 1036
rect 850 1028 853 1031
rect 563 1023 572 1026
rect 494 995 505 998
rect 563 994 572 997
rect 606 993 613 996
rect 490 989 505 992
rect 566 988 572 991
rect 539 975 542 978
rect 566 966 569 988
rect 495 963 569 966
rect 572 963 576 966
rect 610 958 613 993
rect 628 969 632 972
rect 479 955 613 958
rect 479 923 482 955
rect 629 934 632 969
rect 629 931 788 934
rect 348 920 482 923
rect 348 887 351 920
rect 713 892 714 895
rect 348 884 355 887
rect 360 884 361 887
rect -3 876 0 879
rect 354 830 361 833
rect -3 802 0 805
rect 354 784 357 830
rect 354 781 484 784
rect 481 738 484 781
rect 606 762 609 775
rect 568 748 572 751
rect 479 735 484 738
rect 567 742 572 745
rect 630 743 633 746
rect 505 732 509 735
rect 567 734 570 742
rect 563 729 570 734
rect 636 727 643 730
rect 12 718 17 721
rect 636 717 639 727
rect 677 717 680 730
rect 630 714 639 717
rect 606 713 630 714
rect 490 708 507 711
rect 638 686 643 689
rect 701 685 707 688
rect 487 674 490 682
rect 501 680 507 683
rect 628 682 643 683
rect 633 680 643 682
rect 487 671 507 674
rect 640 654 643 664
rect 677 661 680 669
rect 627 651 643 654
rect 363 635 504 638
rect 704 638 707 685
rect 559 635 707 638
rect -3 595 0 598
rect 363 583 366 635
rect 725 588 728 591
rect 363 580 373 583
rect 501 582 502 585
rect 293 526 373 529
rect -3 521 0 524
rect 293 483 296 526
rect 522 492 525 500
rect 293 480 483 483
rect 617 481 620 494
rect 480 457 483 480
rect 579 467 583 470
rect 578 461 583 464
rect 641 462 644 465
rect 508 451 520 454
rect 578 453 581 461
rect 574 448 581 453
rect 647 446 654 449
rect 647 436 650 446
rect 688 436 691 449
rect 641 433 650 436
rect 617 432 641 433
rect 490 427 518 430
rect 649 405 654 408
rect 712 404 718 407
rect 487 393 490 401
rect 513 399 518 402
rect 639 399 654 402
rect 487 390 518 393
rect 487 362 490 390
rect 651 373 654 383
rect 688 380 691 388
rect 715 376 718 404
rect 638 370 654 373
rect 660 373 718 376
rect 317 359 490 362
rect 317 356 320 359
rect 257 353 320 356
rect 660 353 663 373
rect -3 314 0 317
rect -3 237 0 240
rect 257 199 260 353
rect 340 350 663 353
rect 340 296 343 350
rect 715 301 718 304
rect 340 293 363 296
rect 491 295 493 298
rect 257 196 446 199
rect 443 162 446 196
rect 466 190 501 193
rect 706 187 712 190
rect 746 189 749 190
rect 671 184 674 185
rect 706 184 709 187
rect 671 182 709 184
rect 695 181 709 182
rect 443 159 496 162
rect 485 38 488 117
rect 493 91 496 159
rect 620 156 623 165
rect 707 158 712 161
rect 770 157 776 160
rect 620 153 637 156
rect 695 152 712 155
rect 630 147 637 150
rect 613 128 616 139
rect 671 123 674 136
rect 692 131 695 136
rect 692 128 712 131
rect 746 128 749 141
rect 773 125 776 157
rect 716 122 776 125
rect 571 112 579 115
rect 574 106 579 109
rect 637 107 640 110
rect 508 96 516 99
rect 574 98 577 106
rect 570 93 577 98
rect 713 96 719 99
rect 643 91 650 94
rect 643 81 646 91
rect 684 81 687 94
rect 713 81 716 96
rect 753 86 756 99
rect 637 78 646 81
rect 708 78 716 81
rect 613 77 637 78
rect 498 72 514 75
rect 716 55 719 58
rect 785 57 788 931
rect 777 54 788 57
rect 645 50 650 53
rect 708 49 719 52
rect 509 44 514 47
rect 635 44 650 47
rect 485 35 514 38
rect -2 30 1 33
rect 647 18 650 28
rect 684 25 687 33
rect 705 30 719 33
rect 753 30 756 38
rect 634 15 650 18
rect -2 -7 40 -4
rect 45 -7 595 -4
rect 600 -7 614 -4
<< m2contact >>
rect 490 962 495 967
rect 663 940 668 945
rect 663 922 668 927
rect 518 802 523 807
rect 500 732 505 737
rect 633 741 638 746
rect 633 686 638 691
rect 479 680 484 685
rect 496 680 501 685
rect 503 451 508 456
rect 644 460 649 465
rect 644 405 649 410
rect 508 399 513 404
rect 461 189 466 194
rect 501 188 506 193
rect 620 165 625 170
rect 625 145 630 150
rect 711 120 716 125
rect 503 96 508 101
rect 640 105 645 110
rect 492 86 497 91
rect 493 71 498 76
rect 711 55 716 60
rect 640 50 645 55
rect 504 44 509 49
<< metal2 >>
rect 267 1199 296 1202
rect 267 1041 270 1199
rect 295 1120 298 1148
rect 295 1117 372 1120
rect 369 1085 372 1117
rect 369 1082 781 1085
rect 267 1038 484 1041
rect 481 1019 484 1038
rect 479 1014 484 1019
rect 481 979 484 987
rect 481 976 504 979
rect 491 929 494 962
rect 296 926 494 929
rect 296 756 299 926
rect 501 922 504 976
rect 664 927 667 940
rect 303 919 504 922
rect 303 763 306 919
rect 519 776 522 802
rect 549 777 552 865
rect 549 774 596 777
rect 303 760 504 763
rect 296 753 494 756
rect 479 735 484 738
rect 491 728 494 753
rect 501 737 504 760
rect 567 729 623 732
rect 491 725 499 728
rect 12 718 17 721
rect 480 694 483 706
rect 480 691 492 694
rect 480 649 483 680
rect 290 646 483 649
rect 290 475 293 646
rect 489 642 492 691
rect 496 685 499 725
rect 620 648 623 729
rect 635 691 638 741
rect 617 645 623 648
rect 617 644 620 645
rect 297 639 492 642
rect 569 641 620 644
rect 297 482 300 639
rect 569 501 572 641
rect 629 639 632 641
rect 624 637 632 639
rect 576 636 632 637
rect 576 634 627 636
rect 576 524 579 634
rect 576 521 643 524
rect 569 498 623 501
rect 297 479 506 482
rect 290 472 499 475
rect 480 413 483 425
rect 496 420 499 472
rect 503 456 506 479
rect 496 417 511 420
rect 480 410 501 413
rect 498 368 501 410
rect 508 404 511 417
rect 275 365 501 368
rect 275 356 278 365
rect 251 353 278 356
rect 566 363 578 366
rect 251 194 254 353
rect 367 242 372 243
rect 297 239 372 242
rect 297 201 300 239
rect 367 238 372 239
rect 297 198 483 201
rect 251 191 461 194
rect 480 173 483 198
rect 566 189 569 363
rect 620 362 623 498
rect 640 490 643 521
rect 634 487 643 490
rect 646 410 649 460
rect 620 359 641 362
rect 480 75 483 141
rect 503 101 506 188
rect 638 170 641 359
rect 778 185 781 1082
rect 703 182 781 185
rect 625 167 641 170
rect 703 163 706 182
rect 625 98 628 145
rect 574 95 628 98
rect 497 86 508 89
rect 480 72 493 75
rect 505 49 508 86
rect 642 55 645 105
rect 712 60 715 120
<< m123contact >>
rect 97 1270 102 1275
rect 546 1269 551 1274
rect 410 1261 415 1266
rect 244 1181 249 1186
rect 257 1051 262 1056
rect 410 1143 415 1148
rect 539 1036 544 1041
rect 629 1022 634 1027
rect 537 970 542 975
rect 576 963 581 968
rect 355 884 360 889
rect 485 885 490 890
rect 596 772 601 777
rect 551 751 556 756
rect 563 748 568 753
rect 588 651 593 656
rect 597 651 602 656
rect 628 677 633 682
rect 629 641 634 646
rect 504 635 509 640
rect 554 635 559 640
rect 496 582 501 587
rect 609 489 614 494
rect 574 467 579 472
rect 562 461 567 466
rect 599 370 604 375
rect 485 295 491 301
rect 578 362 583 367
rect 629 485 634 490
rect 565 184 570 189
rect 665 182 670 187
rect 702 158 707 163
rect 556 137 561 142
rect 613 123 618 128
rect 566 112 571 117
rect 665 91 670 96
rect 595 15 600 20
rect 40 -8 45 -3
rect 595 -7 600 -2
<< metal3 >>
rect 98 1245 101 1270
rect 246 1115 249 1181
rect 411 1148 414 1261
rect 547 1229 550 1269
rect 443 1159 446 1164
rect 334 1115 337 1135
rect 246 1112 337 1115
rect 411 1091 414 1143
rect 501 1107 504 1112
rect 411 1088 705 1091
rect 258 1046 261 1051
rect 258 1043 347 1046
rect 344 763 347 1043
rect 407 1043 542 1046
rect 407 1030 410 1043
rect 539 1041 542 1043
rect 629 1027 632 1088
rect 539 966 542 970
rect 539 963 576 966
rect 652 967 655 988
rect 581 964 655 967
rect 539 961 542 963
rect 446 958 542 961
rect 446 934 449 958
rect 702 931 705 1088
rect 702 928 735 931
rect 356 784 359 884
rect 486 798 489 885
rect 732 798 735 928
rect 486 795 735 798
rect 356 781 616 784
rect 344 760 567 763
rect 407 753 551 756
rect 407 749 410 753
rect 564 753 567 760
rect 597 656 600 772
rect 449 653 588 656
rect 613 647 616 781
rect 317 644 616 647
rect 629 646 632 677
rect 317 637 320 644
rect 262 634 320 637
rect 509 635 554 638
rect 262 479 265 634
rect 732 630 735 795
rect 497 627 735 630
rect 497 587 500 627
rect 561 552 564 557
rect 561 549 612 552
rect 609 494 612 549
rect 262 476 578 479
rect 575 472 578 476
rect 407 463 562 466
rect 610 375 613 489
rect 446 372 599 375
rect 446 282 449 372
rect 604 372 613 375
rect 629 366 632 485
rect 583 363 632 366
rect 732 348 735 627
rect 486 345 735 348
rect 486 301 489 345
rect 446 279 521 282
rect 368 207 378 210
rect 368 183 371 207
rect 453 149 456 150
rect 453 146 560 149
rect 557 142 560 146
rect 566 117 569 184
rect 41 -3 44 46
rect 614 18 617 123
rect 666 96 669 182
rect 600 15 617 18
rect 596 -2 599 15
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 292 0 1 1105
box -3 -9 349 129
use nor  nor_0
timestamp 1618580541
transform 1 0 505 0 1 1000
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 539 0 1 993
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 572 0 1 999
box 0 -35 34 27
use ffo  ffo_0
timestamp 1618618535
transform 1 0 643 0 -1 1030
box -14 -42 207 91
use sumffo  sumffo_1
timestamp 1618628987
transform 1 0 364 0 -1 927
box -3 -9 349 129
use nand  nand_1
timestamp 1618580231
transform 1 0 572 0 -1 740
box 0 -35 34 27
use inv  inv_1
timestamp 1618579805
transform 1 0 606 0 -1 747
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 683
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 643 0 1 691
box 0 -30 34 39
use inv  inv_2
timestamp 1618579805
transform 1 0 677 0 1 684
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1618628987
transform 1 0 376 0 -1 623
box -3 -9 349 129
use nand  nand_2
timestamp 1618580231
transform 1 0 583 0 -1 459
box 0 -35 34 27
use inv  inv_3
timestamp 1618579805
transform 1 0 617 0 -1 466
box 0 -15 24 33
use cla  cla_1
timestamp 1618627066
transform 1 0 527 0 1 402
box -9 -46 112 95
use nor  nor_2
timestamp 1618580541
transform 1 0 654 0 1 410
box 0 -30 34 39
use inv  inv_4
timestamp 1618579805
transform 1 0 688 0 1 403
box 0 -15 24 33
use sumffo  sumffo_3
timestamp 1618628987
transform 1 0 366 0 -1 336
box -3 -9 349 129
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use nand  nand_3
timestamp 1618580231
transform 1 0 579 0 -1 104
box 0 -35 34 27
use inv  inv_5
timestamp 1618579805
transform 1 0 613 0 -1 111
box 0 -15 24 33
use nand  nand_4
timestamp 1618580231
transform 1 0 637 0 1 158
box 0 -35 34 27
use inv  inv_7
timestamp 1618579805
transform 1 0 671 0 1 151
box 0 -15 24 33
use nand  nand_5
timestamp 1618580231
transform 1 0 712 0 1 163
box 0 -35 34 27
use inv  inv_8
timestamp 1618579805
transform 1 0 746 0 1 156
box 0 -15 24 33
use cla  cla_2
timestamp 1618627066
transform 1 0 523 0 1 47
box -9 -46 112 95
use nor  nor_3
timestamp 1618580541
transform 1 0 650 0 1 55
box 0 -30 34 39
use inv  inv_6
timestamp 1618579805
transform 1 0 684 0 1 48
box 0 -15 24 33
use nor  nor_4
timestamp 1618580541
transform 1 0 719 0 1 60
box 0 -30 34 39
use inv  inv_9
timestamp 1618579805
transform 1 0 753 0 1 53
box 0 -15 24 33
<< labels >>
rlabel metal1 -3 314 -3 317 3 y3in
rlabel metal1 -3 1153 -3 1156 3 cinin
rlabel metal1 -3 1083 -3 1086 3 x1in
rlabel metal1 -3 876 -3 879 3 y1in
rlabel metal1 -3 802 -3 805 3 x2in
rlabel metal1 -3 595 -3 598 3 y2in
rlabel metal1 -3 521 -3 524 3 x3in
rlabel metal1 -3 237 -3 240 3 x4in
rlabel metal1 -2 30 -2 33 3 y4in
rlabel metal1 -3 1252 -3 1255 3 clk
rlabel metal1 71 1271 71 1271 5 vdd!
rlabel metal1 644 1137 644 1140 7 z1o
rlabel metal1 714 892 714 895 7 z2o
rlabel metal1 728 588 728 591 7 z3o
rlabel metal1 718 301 718 304 7 z4o
rlabel metal1 853 1028 853 1031 1 couto
rlabel metal1 19 -6 19 -6 1 gnd!
<< end >>
