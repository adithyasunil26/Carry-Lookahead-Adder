* SPICE3 file created from inv.ext - technology: scmos

.option scale=0.09u

M1000 op in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=30 ps=22
M1001 op in vdd w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=60 ps=34
C0 gnd op 0.10fF
C1 gnd in 0.05fF
C2 op vdd 0.15fF
C3 op in 0.04fF
C4 vdd in 0.02fF
C5 op w_0_6# 0.03fF
C6 vdd w_0_6# 0.06fF
C7 in w_0_6# 0.06fF
C8 gnd Gnd 0.09fF
C9 op Gnd 0.05fF
C10 vdd Gnd 0.03fF
C11 in Gnd 0.14fF
C12 w_0_6# Gnd 0.58fF
