* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 vdd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 vdd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 s1 cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op s1 sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op s1 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 s1 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 vdd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 sumffo_2/xor_0/op ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_2/xor_0/op sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 s2 nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op s2 sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op s2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 s2 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 vdd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 s4 ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op s4 sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op s4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 s4 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 vdd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in vdd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 vdd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in vdd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in vdd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 vdd y2in cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 cla_1/g0 x2in vdd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_1/g0 y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 vdd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in vdd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in vdd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 vdd y3in cla_2/g0 ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1196 cla_2/g0 x3in vdd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_2/g0 y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 vdd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in vdd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in vdd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 vdd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in vdd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 vdd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in vdd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in vdd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C1 cla_0/nor_1/w_0_0# vdd 0.31fF
C2 cin sumffo_3/xor_0/a_10_10# 0.04fF
C3 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C4 x1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C5 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/op 0.02fF
C6 cla_0/g0 cin 0.08fF
C7 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C8 cla_1/g0 gnd 0.28fF
C9 cla_1/g0 cla_1/p0 0.07fF
C10 nand_2/b cla_0/n 0.06fF
C11 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C12 cla_2/g1 gnd 0.30fF
C13 vdd ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C14 y3in ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C15 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C16 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C17 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C18 vdd sumffo_3/xor_0/a_10_10# 0.93fF
C19 cla_0/g0 vdd 0.54fF
C20 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C21 ffipg_2/k cla_0/n 0.06fF
C22 nand_2/b inv_3/w_0_6# 0.06fF
C23 cla_2/p0 y3in 0.03fF
C24 vdd ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C25 cla_0/inv_0/in vdd 0.05fF
C26 cla_2/nor_1/w_0_0# vdd 0.31fF
C27 cin sumffo_1/xor_0/inv_1/op 0.04fF
C28 y3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C29 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.17fF
C30 inv_3/in nor_2/b 0.04fF
C31 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C32 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C33 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C34 vdd sumffo_3/xor_0/inv_0/op 0.15fF
C35 ffipg_3/pggen_0/xor_0/inv_0/op x4in 0.27fF
C36 cla_0/nand_0/w_0_0# vdd 0.10fF
C37 inv_9/in cout 0.04fF
C38 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C39 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C40 inv_8/w_0_6# inv_8/in 0.10fF
C41 vdd ffipg_3/pggen_0/xor_0/inv_1/op 0.15fF
C42 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C43 vdd sumffo_1/xor_0/inv_1/op 0.15fF
C44 vdd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C45 cla_1/l vdd 0.22fF
C46 cin sumffo_0/xor_0/inv_0/op 0.20fF
C47 gnd inv_7/in 0.13fF
C48 inv_7/w_0_6# inv_7/in 0.10fF
C49 y2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C50 gnd inv_2/in 0.17fF
C51 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C52 cla_0/g0 y1in 0.13fF
C53 cin sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C54 inv_2/w_0_6# inv_2/in 0.10fF
C55 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C56 vdd nor_4/a 0.19fF
C57 vdd sumffo_0/xor_0/inv_0/op 0.15fF
C58 ffipg_2/pggen_0/xor_0/inv_1/op y3in 0.22fF
C59 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C60 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C61 inv_1/op inv_1/in 0.04fF
C62 gnd s4 0.14fF
C63 cla_2/g0 cla_2/inv_0/in 0.16fF
C64 vdd sumffo_0/xor_0/inv_1/w_0_6# 0.07fF
C65 gnd y4in 1.66fF
C66 cla_1/l cla_0/n 0.07fF
C67 ffipg_1/k x2in 0.46fF
C68 gnd cout 0.10fF
C69 y1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C70 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C71 cla_0/l cla_2/g0 0.05fF
C72 cla_2/p1 cla_2/inv_0/in 0.02fF
C73 vdd nor_3/b 0.23fF
C74 vdd cla_2/inv_0/op 0.17fF
C75 x1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C76 gnd ffipg_3/k 0.31fF
C77 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C78 cla_1/l inv_3/w_0_6# 0.06fF
C79 cla_0/l cla_0/inv_0/w_0_6# 0.00fF
C80 vdd nor_1/w_0_0# 0.17fF
C81 gnd inv_4/in 0.24fF
C82 nand_2/b inv_3/in 0.13fF
C83 vdd cla_2/n 0.28fF
C84 gnd x2in 0.31fF
C85 ffipg_0/k x1in 0.46fF
C86 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C87 gnd x3in 0.31fF
C88 cla_1/p0 x2in 0.22fF
C89 vdd inv_9/in 0.09fF
C90 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C91 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C92 ffipg_3/pggen_0/xor_0/w_n3_4# x4in 0.06fF
C93 cla_2/l nor_3/b 0.10fF
C94 cla_2/g0 cla_2/p0 0.08fF
C95 cla_0/inv_0/op vdd 0.17fF
C96 cin ffipg_1/k 0.06fF
C97 cla_2/g0 ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C98 gnd x1in 0.22fF
C99 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C100 cla_1/nand_0/w_0_0# gnd 0.01fF
C101 cla_2/g1 y4in 0.13fF
C102 vdd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C103 inv_7/op inv_8/w_0_6# 0.06fF
C104 cla_1/inv_0/in gnd 0.30fF
C105 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C106 cla_0/l nand_2/b 0.08fF
C107 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C108 sumffo_1/xor_0/a_10_10# s2 0.45fF
C109 cla_2/p0 cla_2/p1 0.24fF
C110 cin ffipg_0/k 0.19fF
C111 vdd ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C112 nor_1/w_0_0# cla_0/n 0.06fF
C113 vdd ffipg_1/k 0.36fF
C114 cla_1/inv_0/op gnd 0.10fF
C115 cla_0/l ffipg_2/k 0.04fF
C116 cla_1/nor_0/w_0_0# vdd 0.31fF
C117 cin gnd 0.74fF
C118 sumffo_0/xor_0/w_n3_4# s1 0.02fF
C119 vdd ffipg_0/k 0.33fF
C120 cin inv_2/w_0_6# 0.06fF
C121 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C122 nor_2/w_0_0# inv_4/in 0.11fF
C123 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C124 nor_1/w_0_0# nor_1/b 0.06fF
C125 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C126 vdd gnd 3.74fF
C127 vdd inv_7/w_0_6# 0.15fF
C128 nor_0/w_0_0# nor_0/a 0.06fF
C129 cla_1/p0 vdd 0.43fF
C130 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.02fF
C131 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C132 cla_1/g0 cla_1/inv_0/in 0.16fF
C133 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C134 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C135 vdd inv_2/w_0_6# 0.15fF
C136 ffipg_2/pggen_0/xor_0/w_n3_4# x3in 0.06fF
C137 cla_2/p0 ffipg_2/k 0.05fF
C138 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C139 vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C140 cin sumffo_1/xor_0/a_38_n43# 0.01fF
C141 y1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C142 x1in ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C143 cla_0/l cla_0/inv_0/in 0.14fF
C144 cla_2/l gnd 0.24fF
C145 cla_2/l inv_7/w_0_6# 0.06fF
C146 y4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C147 nor_3/w_0_0# nor_3/b 0.06fF
C148 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C149 cin sumffo_1/xor_0/w_n3_4# 0.00fF
C150 ffipg_0/k y1in 0.07fF
C151 ffipg_0/pggen_0/nand_0/w_0_0# x1in 0.06fF
C152 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C153 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C154 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C155 cla_0/l cla_0/nand_0/w_0_0# 0.00fF
C156 cla_2/p1 x4in 0.22fF
C157 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C158 y2in ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C159 gnd cla_0/n 0.61fF
C160 vdd ffipg_1/pggen_0/nand_0/a_13_n26# 0.01fF
C161 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C162 cla_1/g0 vdd 0.55fF
C163 nor_3/w_0_0# cla_2/n 0.06fF
C164 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C165 cla_2/g1 vdd 0.35fF
C166 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C167 cin sumffo_2/xor_0/a_10_10# 0.04fF
C168 gnd y1in 1.64fF
C169 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C170 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C171 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.21fF
C172 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C173 x2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C174 y2in ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C175 vdd sumffo_1/xor_0/w_n3_4# 0.12fF
C176 gnd inv_3/w_0_6# 0.02fF
C177 ffipg_3/k y4in 0.07fF
C178 vdd nor_2/w_0_0# 0.17fF
C179 cin sumffo_1/xor_0/inv_0/op 0.06fF
C180 nor_0/a cinbar 0.32fF
C181 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C182 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C183 y2in ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C184 vdd ffipg_0/pggen_0/xor_0/inv_0/op 0.15fF
C185 vdd sumffo_2/xor_0/a_10_10# 0.93fF
C186 vdd ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C187 gnd nor_1/b 0.10fF
C188 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C189 inv_2/w_0_6# nor_1/b 0.03fF
C190 vdd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C191 vdd sumffo_1/xor_0/inv_0/op 0.15fF
C192 cin inv_2/in 0.13fF
C193 cla_1/g0 cla_0/n 0.13fF
C194 cla_1/l cla_2/p0 0.02fF
C195 cla_1/inv_0/w_0_6# vdd 0.06fF
C196 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C197 cla_2/g0 y3in 0.13fF
C198 inv_0/in nor_0/a 0.02fF
C199 vdd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C200 sumffo_0/xor_0/inv_0/w_0_6# ffipg_0/k 0.06fF
C201 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C202 vdd inv_7/in 0.30fF
C203 nor_0/w_0_0# cinbar 0.06fF
C204 cin s4 0.16fF
C205 vdd inv_2/in 0.30fF
C206 nor_4/a nor_4/w_0_0# 0.07fF
C207 sumffo_0/xor_0/inv_0/w_0_6# gnd 0.02fF
C208 vdd ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C209 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C210 inv_5/w_0_6# inv_5/in 0.10fF
C211 y1in ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C212 gnd inv_4/op 0.32fF
C213 vdd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C214 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C215 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C216 y4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C217 inv_6/in nor_3/b 0.16fF
C218 sumffo_3/xor_0/inv_1/op s4 0.52fF
C219 nor_0/w_0_0# inv_0/in 0.11fF
C220 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C221 ffipg_0/pggen_0/nand_0/w_0_0# y1in 0.06fF
C222 gnd sumffo_2/xor_0/op 0.14fF
C223 nor_0/w_0_0# inv_0/op 0.10fF
C224 cla_0/l cla_0/inv_0/op 0.21fF
C225 cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C226 vdd y4in 0.10fF
C227 vdd cout 0.15fF
C228 vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C229 inv_6/in cla_2/n 0.02fF
C230 inv_8/w_0_6# nor_4/a 0.03fF
C231 inv_1/op ffipg_2/k 0.09fF
C232 s1 sumffo_0/xor_0/inv_0/op 0.06fF
C233 vdd ffipg_3/k 0.35fF
C234 ffipg_3/pggen_0/xor_0/inv_1/op x4in 0.06fF
C235 sumffo_2/xor_0/inv_0/op gnd 0.17fF
C236 gnd inv_3/in 0.17fF
C237 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C238 vdd inv_4/in 0.09fF
C239 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C240 nor_4/b nor_4/a 0.42fF
C241 cin sumffo_0/xor_0/a_10_10# 0.12fF
C242 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C243 ffipg_2/k y3in 0.07fF
C244 inv_9/in nor_4/w_0_0# 0.11fF
C245 vdd x2in 0.93fF
C246 vdd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C247 vdd x3in 0.93fF
C248 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/inv_0/op 0.08fF
C249 nor_0/w_0_0# nand_2/b 0.04fF
C250 inv_2/in nor_1/b 0.04fF
C251 cla_2/inv_0/in gnd 0.30fF
C252 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C253 vdd x1in 0.97fF
C254 inv_4/op nor_2/w_0_0# 0.03fF
C255 vdd sumffo_0/xor_0/a_10_10# 0.93fF
C256 cla_1/nand_0/w_0_0# vdd 0.10fF
C257 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C258 cla_1/inv_0/in vdd 0.05fF
C259 cla_0/l inv_7/w_0_6# 0.06fF
C260 cla_0/l gnd 0.98fF
C261 cla_0/l cla_1/p0 0.02fF
C262 ffipg_3/k cla_0/n 0.06fF
C263 inv_0/in cinbar 0.16fF
C264 cla_0/l inv_2/w_0_6# 0.06fF
C265 cla_0/g0 nor_0/a 0.40fF
C266 ffipg_1/k y2in 0.07fF
C267 nor_2/b cla_1/n 0.39fF
C268 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/op 0.45fF
C269 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C270 cla_1/inv_0/op vdd 0.17fF
C271 cla_0/nand_0/a_13_n26# gnd 0.00fF
C272 gnd inv_6/in 0.24fF
C273 vdd cin 2.44fF
C274 cin sumffo_3/xor_0/inv_1/op 0.04fF
C275 nor_4/b inv_9/in 0.16fF
C276 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C277 vdd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C278 ffipg_2/pggen_0/xor_0/inv_0/op x3in 0.27fF
C279 cla_2/g1 cla_2/inv_0/in 0.04fF
C280 cla_2/p0 gnd 0.68fF
C281 vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C282 cla_2/g0 cla_2/p1 0.30fF
C283 cla_1/p0 cla_2/p0 0.24fF
C284 inv_1/in nor_1/w_0_0# 0.11fF
C285 inv_0/op inv_0/in 0.04fF
C286 gnd y2in 1.68fF
C287 x1in y1in 0.73fF
C288 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C289 nor_0/w_0_0# cla_0/g0 0.06fF
C290 cla_0/l cla_1/g0 0.12fF
C291 vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C292 cla_1/p0 y2in 0.03fF
C293 vdd sumffo_3/xor_0/inv_1/op 0.15fF
C294 cla_2/g0 cla_1/n 0.13fF
C295 cla_1/inv_0/op cla_0/n 0.06fF
C296 inv_8/in nor_4/a 0.04fF
C297 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C298 vdd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C299 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C300 cla_2/l vdd 0.38fF
C301 x2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C302 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C303 cla_1/nor_1/w_0_0# vdd 0.31fF
C304 gnd s1 0.14fF
C305 cin sumffo_0/xor_0/inv_1/op 0.22fF
C306 vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C307 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C308 cla_1/g0 cla_2/p0 0.36fF
C309 ffipg_3/k inv_4/op 0.09fF
C310 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C311 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C312 vdd cla_0/n 0.56fF
C313 gnd nor_4/b 0.10fF
C314 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.24fF
C315 x2in ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C316 cla_1/g0 y2in 0.13fF
C317 vdd y1in 0.15fF
C318 inv_4/op inv_4/in 0.04fF
C319 vdd sumffo_0/xor_0/inv_1/op 0.15fF
C320 vdd ffipg_2/pggen_0/xor_0/inv_0/op 0.15fF
C321 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C322 inv_1/op nor_1/w_0_0# 0.03fF
C323 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C324 cla_0/l inv_7/in 0.13fF
C325 vdd inv_3/w_0_6# 0.15fF
C326 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C327 gnd x4in 0.31fF
C328 cla_2/l cla_0/n 0.32fF
C329 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C330 y1in ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C331 vdd nor_1/b 0.25fF
C332 gnd inv_1/in 0.24fF
C333 inv_5/w_0_6# nor_3/b 0.17fF
C334 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.21fF
C335 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C336 y1in ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C337 vdd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C338 cla_2/g0 cla_2/nor_1/w_0_0# 0.06fF
C339 sumffo_3/xor_0/w_n3_4# s4 0.02fF
C340 inv_0/op cla_0/g0 0.32fF
C341 ffipg_2/k nand_2/b 0.06fF
C342 inv_3/w_0_6# cla_0/n 0.16fF
C343 y3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C344 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C345 ffipg_1/k nor_0/a 0.06fF
C346 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C347 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C348 vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C349 cla_0/l ffipg_3/k 0.04fF
C350 sumffo_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C351 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C352 vdd nor_3/w_0_0# 0.14fF
C353 cin sumffo_2/xor_0/op 0.27fF
C354 nor_1/b cla_0/n 0.36fF
C355 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C356 y2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C357 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C358 vdd inv_4/op 0.26fF
C359 cla_2/nand_0/w_0_0# gnd 0.08fF
C360 ffipg_0/k nor_0/a 0.05fF
C361 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C362 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C363 gnd inv_1/op 0.32fF
C364 gnd inv_8/in 0.13fF
C365 cout nor_4/w_0_0# 0.03fF
C366 sumffo_2/xor_0/inv_0/op cin 0.06fF
C367 gnd nor_0/a 0.23fF
C368 cla_1/p0 nor_0/a 0.24fF
C369 sumffo_1/xor_0/inv_1/op s2 0.52fF
C370 cla_0/l cla_1/nand_0/w_0_0# 0.01fF
C371 cla_0/g0 nand_2/b 0.13fF
C372 gnd y3in 1.68fF
C373 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C374 cla_2/p0 ffipg_3/k 0.06fF
C375 vdd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C376 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C377 sumffo_2/xor_0/inv_0/op vdd 0.15fF
C378 vdd inv_3/in 0.30fF
C379 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C380 gnd inv_5/w_0_6# 0.26fF
C381 cla_0/l cla_1/inv_0/op 0.05fF
C382 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# y3in 0.23fF
C383 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C384 cla_2/p0 x3in 0.22fF
C385 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C386 cin sumffo_3/xor_0/a_38_n43# 0.01fF
C387 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C388 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C389 cla_0/l cin 0.33fF
C390 x3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C391 x2in y2in 0.73fF
C392 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C393 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C394 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C395 vdd cla_2/inv_0/in 0.05fF
C396 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C397 cla_1/l nand_2/b 0.31fF
C398 inv_5/in nor_3/b 0.04fF
C399 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C400 cla_1/inv_0/in cla_2/p0 0.02fF
C401 cla_0/l vdd 0.53fF
C402 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C403 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C404 vdd cla_2/inv_0/w_0_6# 0.06fF
C405 cin sumffo_1/xor_0/a_10_10# 0.04fF
C406 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C407 cla_0/g0 cla_0/inv_0/in 0.16fF
C408 y4in x4in 0.73fF
C409 vdd inv_6/in 0.09fF
C410 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C411 s1 sumffo_0/xor_0/a_10_10# 0.45fF
C412 inv_3/w_0_6# inv_3/in 0.10fF
C413 vdd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C414 cla_0/l cla_2/l 0.37fF
C415 ffipg_2/pggen_0/xor_0/inv_1/op x3in 0.06fF
C416 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C417 vdd sumffo_1/xor_0/a_10_10# 0.93fF
C418 ffipg_0/k cinbar 0.06fF
C419 ffipg_3/pggen_0/xor_0/inv_0/op y4in 0.20fF
C420 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C421 gnd nor_2/b 0.10fF
C422 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C423 ffipg_3/k x4in 0.46fF
C424 vdd nor_4/w_0_0# 0.15fF
C425 cla_2/p0 vdd 0.43fF
C426 cin sumffo_2/xor_0/inv_1/op 0.04fF
C427 vdd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C428 y2in ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C429 inv_7/op gnd 0.10fF
C430 inv_7/op inv_7/w_0_6# 0.03fF
C431 cla_0/l cla_0/n 0.05fF
C432 vdd y2in 0.15fF
C433 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C434 ffipg_3/k sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C435 cin inv_8/w_0_6# 0.06fF
C436 cla_0/l inv_3/w_0_6# 0.00fF
C437 vdd sumffo_2/xor_0/inv_1/op 0.15fF
C438 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C439 cla_2/l cla_2/p0 0.16fF
C440 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C441 cla_0/inv_0/op nand_2/b 0.09fF
C442 cla_2/g0 gnd 0.27fF
C443 vdd inv_8/w_0_6# 0.15fF
C444 gnd inv_5/in 0.19fF
C445 gnd inv_0/in 0.24fF
C446 ffipg_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C447 inv_0/op gnd 0.10fF
C448 vdd nor_4/b 0.15fF
C449 cla_2/p1 gnd 0.68fF
C450 vdd ffipg_2/pggen_0/xor_0/inv_1/op 0.15fF
C451 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C452 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C453 nor_2/b nor_2/w_0_0# 0.06fF
C454 gnd s2 0.14fF
C455 nand_2/b ffipg_1/k 0.15fF
C456 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C457 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C458 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op 0.06fF
C459 gnd cla_1/n 0.23fF
C460 vdd x4in 0.93fF
C461 vdd inv_1/in 0.09fF
C462 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# x4in 0.06fF
C463 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C464 cla_1/g0 cla_2/g0 0.35fF
C465 vdd ffipg_2/pggen_0/nand_0/a_13_n26# 0.01fF
C466 cla_2/g0 cla_2/g1 0.26fF
C467 cla_2/nor_0/w_0_0# vdd 0.31fF
C468 s1 sumffo_0/xor_0/inv_1/op 0.52fF
C469 gnd nand_2/b 0.83fF
C470 vdd ffipg_3/pggen_0/xor_0/inv_0/op 0.15fF
C471 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C472 y3in x3in 0.73fF
C473 vdd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C474 nand_2/b inv_2/w_0_6# 0.03fF
C475 ffipg_3/pggen_0/xor_0/w_n3_4# y4in 0.06fF
C476 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C477 nor_0/a x1in 0.22fF
C478 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C479 y2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C480 nor_3/w_0_0# inv_6/in 0.11fF
C481 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C482 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C483 cla_2/g1 cla_2/p1 0.00fF
C484 gnd ffipg_2/k 0.29fF
C485 cla_1/p0 ffipg_2/k 0.06fF
C486 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C487 inv_7/op inv_7/in 0.04fF
C488 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C489 vdd ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C490 cla_1/nand_0/a_13_n26# gnd 0.01fF
C491 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C492 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C493 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C494 sumffo_1/xor_0/w_n3_4# s2 0.02fF
C495 cla_0/g0 ffipg_1/k 0.06fF
C496 cin inv_8/in 0.13fF
C497 x2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C498 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C499 cla_0/l inv_3/in 0.22fF
C500 inv_1/in cla_0/n 0.02fF
C501 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C502 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# y4in 0.23fF
C503 nor_2/w_0_0# cla_1/n 0.06fF
C504 cla_2/nand_0/w_0_0# vdd 0.10fF
C505 cla_1/g0 nand_2/b 0.06fF
C506 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.24fF
C507 vdd inv_1/op 0.26fF
C508 vdd inv_8/in 0.30fF
C509 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C510 nor_4/a inv_9/in 0.02fF
C511 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C512 sumffo_1/xor_0/inv_0/op s2 0.06fF
C513 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C514 vdd nor_0/a 0.35fF
C515 cla_0/g0 gnd 0.70fF
C516 cla_0/g0 cla_1/p0 0.38fF
C517 cla_1/g0 ffipg_2/k 0.06fF
C518 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.21fF
C519 cla_0/inv_0/in gnd 0.30fF
C520 inv_1/in nor_1/b 0.16fF
C521 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C522 cla_0/inv_0/in cla_1/p0 0.02fF
C523 vdd y3in 0.15fF
C524 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C525 y1in ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C526 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C527 nor_2/b inv_4/in 0.16fF
C528 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C529 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C530 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op 0.52fF
C531 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C532 nor_0/w_0_0# cin 0.16fF
C533 cla_0/nand_0/w_0_0# gnd 0.01fF
C534 y4in ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C535 nor_3/w_0_0# nor_4/b 0.03fF
C536 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C537 cla_0/nor_0/w_0_0# vdd 0.31fF
C538 cla_2/n nor_3/b 0.41fF
C539 vdd inv_5/w_0_6# 0.15fF
C540 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C541 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C542 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C543 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C544 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C545 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C546 nor_0/w_0_0# vdd 0.46fF
C547 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C548 cla_1/l gnd 0.18fF
C549 vdd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C550 cla_1/p0 cla_1/l 0.16fF
C551 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C552 cin sumffo_2/xor_0/a_38_n43# 0.01fF
C553 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C554 cla_2/g0 ffipg_3/k 0.06fF
C555 cla_2/p1 y4in 0.03fF
C556 vdd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C557 cla_0/g0 cla_1/g0 0.14fF
C558 nand_2/b inv_2/in 0.34fF
C559 nor_0/a y1in 0.03fF
C560 cla_1/g0 cla_0/inv_0/in 0.04fF
C561 cla_2/l inv_5/w_0_6# 0.08fF
C562 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C563 cin sumffo_2/xor_0/w_n3_4# 0.00fF
C564 gnd nor_4/a 0.21fF
C565 sumffo_2/xor_0/inv_1/w_0_6# ffipg_2/k 0.23fF
C566 gnd sumffo_0/xor_0/inv_0/op 0.21fF
C567 cla_2/p1 ffipg_3/k 0.05fF
C568 y3in ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C569 cla_0/nand_0/w_0_0# cla_1/g0 0.06fF
C570 cla_0/n inv_5/w_0_6# 0.06fF
C571 inv_7/op cin 0.31fF
C572 vdd ffipg_0/pggen_0/nand_0/a_13_n26# 0.01fF
C573 vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C574 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C575 cla_2/g0 cla_1/nand_0/w_0_0# 0.06fF
C576 vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C577 cla_2/g0 cla_1/inv_0/in 0.04fF
C578 inv_4/in cla_1/n 0.02fF
C579 vdd nor_2/b 0.21fF
C580 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C581 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C582 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C583 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C584 gnd nor_3/b 0.10fF
C585 cla_2/inv_0/op gnd 0.10fF
C586 inv_7/op vdd 0.17fF
C587 cla_2/g0 cla_1/inv_0/op 0.35fF
C588 vdd cinbar 0.16fF
C589 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C590 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C591 sumffo_0/xor_0/w_n3_4# cin 0.06fF
C592 gnd cla_2/n 0.32fF
C593 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C594 cin inv_0/in 0.07fF
C595 gnd inv_9/in 0.24fF
C596 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C597 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C598 vdd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C599 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# x3in 0.06fF
C600 cla_0/inv_0/op gnd 0.10fF
C601 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C602 inv_6/in nor_4/b 0.04fF
C603 cla_2/g0 vdd 0.55fF
C604 sumffo_3/xor_0/a_10_10# s4 0.45fF
C605 vdd sumffo_0/xor_0/w_n3_4# 0.12fF
C606 vdd inv_5/in 0.30fF
C607 cin s2 0.27fF
C608 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C609 x1in ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C610 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C611 ffipg_2/k x3in 0.46fF
C612 vdd inv_0/in 0.07fF
C613 nor_4/b nor_4/w_0_0# 0.06fF
C614 inv_0/op vdd 0.17fF
C615 cla_2/nand_0/a_13_n26# gnd 0.01fF
C616 cla_0/inv_0/w_0_6# vdd 0.06fF
C617 sumffo_3/xor_0/inv_0/op s4 0.06fF
C618 cla_2/p1 vdd 0.31fF
C619 cla_2/g1 cla_2/inv_0/op 0.35fF
C620 inv_3/w_0_6# nor_2/b 0.03fF
C621 gnd ffipg_1/k 0.39fF
C622 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C623 cla_1/p0 ffipg_1/k 0.05fF
C624 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C625 cla_2/l inv_5/in 0.05fF
C626 cla_2/g0 cla_1/nor_1/w_0_0# 0.02fF
C627 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C628 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C629 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C630 cla_2/g1 cla_2/n 0.13fF
C631 vdd cla_1/n 0.28fF
C632 cin nand_2/b 0.04fF
C633 gnd ffipg_0/k 0.41fF
C634 x2in ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C635 vdd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C636 ffipg_3/pggen_0/xor_0/inv_1/op y4in 0.22fF
C637 cla_0/inv_0/op cla_1/g0 0.35fF
C638 cla_2/g0 cla_0/n 0.06fF
C639 cla_2/l cla_2/p1 0.02fF
C640 ffipg_3/k sumffo_3/xor_0/inv_0/op 0.20fF
C641 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C642 cla_0/n inv_5/in 0.13fF
C643 x2in ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C644 cla_1/p0 gnd 0.68fF
C645 vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C646 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C647 vdd nand_2/b 0.92fF
C648 vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C649 gnd inv_2/w_0_6# 0.02fF
C650 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C651 vdd ffipg_2/k 0.35fF
C652 cla_0/l nor_0/a 0.16fF
C653 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C654 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C655 s3 Gnd 0.00fF **FLOATING
C656 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C657 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C658 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C659 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C660 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C661 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C662 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C663 y4in Gnd 2.72fF
C664 x4in Gnd 2.80fF
C665 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C666 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C667 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C668 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C669 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C670 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C671 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C672 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C673 y3in Gnd 2.72fF
C674 x3in Gnd 2.80fF
C675 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C676 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C677 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C678 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C679 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C680 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C681 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C682 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C683 y2in Gnd 2.72fF
C684 x2in Gnd 2.80fF
C685 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C686 cout Gnd 0.19fF
C687 inv_9/in Gnd 0.23fF
C688 nor_4/w_0_0# Gnd 1.81fF
C689 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C690 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C691 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C692 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C693 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C694 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C695 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C696 y1in Gnd 2.72fF
C697 x1in Gnd 2.80fF
C698 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C699 nor_4/a Gnd 0.59fF
C700 inv_8/in Gnd 0.22fF
C701 inv_8/w_0_6# Gnd 1.40fF
C702 inv_7/in Gnd 0.22fF
C703 inv_7/w_0_6# Gnd 1.40fF
C704 nor_4/b Gnd 0.32fF
C705 nor_3/b Gnd 0.77fF
C706 inv_5/in Gnd 0.22fF
C707 inv_5/w_0_6# Gnd 1.40fF
C708 cla_2/n Gnd 0.36fF
C709 inv_6/in Gnd 0.23fF
C710 nor_3/w_0_0# Gnd 1.81fF
C711 cla_1/n Gnd 0.36fF
C712 inv_4/in Gnd 0.23fF
C713 nor_2/w_0_0# Gnd 1.81fF
C714 cla_0/n Gnd 1.34fF
C715 nor_2/b Gnd 0.70fF
C716 inv_3/in Gnd 0.22fF
C717 inv_3/w_0_6# Gnd 1.40fF
C718 cinbar Gnd 1.15fF
C719 nor_0/a Gnd 1.99fF
C720 nor_1/b Gnd 0.63fF
C721 inv_2/in Gnd 0.22fF
C722 inv_2/w_0_6# Gnd 1.40fF
C723 inv_1/in Gnd 0.23fF
C724 nor_1/w_0_0# Gnd 1.81fF
C725 inv_0/in Gnd 0.23fF
C726 s4 Gnd 0.07fF
C727 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C728 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C729 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C730 ffipg_3/k Gnd 2.89fF
C731 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C732 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C733 inv_4/op Gnd 1.37fF
C734 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C735 s2 Gnd 0.07fF
C736 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C737 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C738 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C739 nand_2/b Gnd 2.99fF
C740 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C741 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C742 ffipg_1/k Gnd 3.04fF
C743 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C744 sumffo_2/xor_0/op Gnd 0.07fF
C745 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C746 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C747 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C748 vdd Gnd 7.86fF
C749 ffipg_2/k Gnd 3.13fF
C750 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C751 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C752 inv_1/op Gnd 1.37fF
C753 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C754 s1 Gnd 0.05fF
C755 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C756 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C757 gnd Gnd 22.85fF
C758 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C759 cin Gnd 6.77fF
C760 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C761 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C762 ffipg_0/k Gnd 2.68fF
C763 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C764 cla_2/p1 Gnd 1.09fF
C765 cla_2/nor_1/w_0_0# Gnd 1.23fF
C766 cla_2/nor_0/w_0_0# Gnd 1.23fF
C767 cla_2/inv_0/in Gnd 0.27fF
C768 cla_2/inv_0/w_0_6# Gnd 0.58fF
C769 cla_2/g1 Gnd 0.59fF
C770 cla_2/inv_0/op Gnd 0.26fF
C771 cla_2/nand_0/w_0_0# Gnd 0.82fF
C772 cla_2/p0 Gnd 0.83fF
C773 cla_1/nor_1/w_0_0# Gnd 1.23fF
C774 cla_1/l Gnd 0.30fF
C775 cla_1/nor_0/w_0_0# Gnd 1.23fF
C776 cla_1/inv_0/in Gnd 0.27fF
C777 cla_1/inv_0/w_0_6# Gnd 0.58fF
C778 cla_2/g0 Gnd 1.58fF
C779 cla_1/inv_0/op Gnd 0.26fF
C780 cla_1/nand_0/w_0_0# Gnd 0.82fF
C781 inv_7/op Gnd 0.26fF
C782 cla_1/p0 Gnd 2.69fF
C783 cla_0/nor_1/w_0_0# Gnd 1.23fF
C784 cla_0/nor_0/w_0_0# Gnd 1.23fF
C785 cla_0/inv_0/in Gnd 0.27fF
C786 cla_0/inv_0/w_0_6# Gnd 0.58fF
C787 cla_1/g0 Gnd 1.59fF
C788 cla_0/inv_0/op Gnd 0.26fF
C789 cla_0/nand_0/w_0_0# Gnd 0.82fF
C790 cla_2/l Gnd 0.25fF
C791 cla_0/g0 Gnd 1.32fF
C792 inv_0/op Gnd 0.23fF
C793 nor_0/w_0_0# Gnd 2.63fF
