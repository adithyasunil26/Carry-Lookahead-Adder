* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 vdd a_35_n5# a_30_8# w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=144 ps=60
M1005 a_7_8# a vdd w_n6_2# pfet w=24 l=2
+  ad=144 pd=60 as=0 ps=0
M1006 a_30_n33# a_27_n20# op Gnd nfet w=12 l=2
+  ad=72 pd=36 as=156 ps=50
M1007 op a_12_3# a_7_8# w_n6_2# pfet w=24 l=2
+  ad=312 pd=74 as=0 ps=0
M1008 gnd a_35_n5# a_30_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_7_n33# a gnd Gnd nfet w=12 l=2
+  ad=72 pd=36 as=0 ps=0
M1010 op b a_7_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_30_8# b op w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 m2_n15_10# inv_0/op 0.02fF
C1 m1_35_n5# op 0.07fF
C2 w_n6_2# inv_1/op 0.09fF
C3 m2_35_n5# m1_35_n5# 0.01fF
C4 inv_0/op vdd 0.15fF
C5 w_n6_2# b 0.16fF
C6 a_35_n5# op 0.06fF
C7 m2_35_n5# inv_0/op 0.02fF
C8 gnd inv_1/op 0.12fF
C9 m2_35_n5# m2_n15_10# 0.02fF
C10 m2_35_n5# a_35_n5# 0.00fF
C11 inv_0/op a 0.08fF
C12 gnd b 0.13fF
C13 a_27_n20# inv_1/op 0.03fF
C14 m2_35_n5# op 0.01fF
C15 vdd a 0.03fF
C16 inv_1/op b 0.44fF
C17 m2_35_n5# a 0.04fF
C18 a_12_3# a 0.03fF
C19 inv_1/op inv_1/w_0_6# 0.04fF
C20 a_35_n5# w_n6_2# 0.06fF
C21 b inv_1/w_0_6# 0.08fF
C22 w_n6_2# vdd 0.09fF
C23 gnd inv_0/op 0.12fF
C24 w_n6_2# op 0.02fF
C25 w_n6_2# a 0.06fF
C26 a_12_3# w_n6_2# 0.08fF
C27 a_27_n20# a_35_n5# 0.04fF
C28 inv_0/op inv_0/w_0_6# 0.04fF
C29 inv_1/op vdd 0.15fF
C30 gnd a 0.42fF
C31 a_35_n5# b 0.04fF
C32 inv_1/op op 0.20fF
C33 m2_35_n5# inv_1/op 0.25fF
C34 vdd inv_0/w_0_6# 0.06fF
C35 b vdd 0.03fF
C36 inv_1/op a 0.15fF
C37 op b 0.22fF
C38 m2_35_n5# b 0.05fF
C39 a_12_3# inv_1/op 0.07fF
C40 a inv_0/w_0_6# 0.08fF
C41 b a 0.11fF
C42 inv_1/w_0_6# vdd 0.06fF
C43 a_35_n5# m1_35_n5# 0.08fF
C44 m2_35_n5# Gnd 0.16fF **FLOATING
C45 m2_n15_10# Gnd 0.09fF **FLOATING
C46 m1_35_n5# Gnd 0.02fF **FLOATING
C47 a_27_n20# Gnd 0.09fF
C48 op Gnd 0.14fF
C49 a_35_n5# Gnd 0.18fF
C50 w_n6_2# Gnd 1.99fF
C51 gnd Gnd 0.39fF
C52 inv_1/op Gnd 0.38fF
C53 b Gnd 1.41fF
C54 inv_1/w_0_6# Gnd 0.58fF
C55 inv_0/op Gnd 0.08fF
C56 vdd Gnd 0.23fF
C57 a Gnd 1.10fF
C58 inv_0/w_0_6# Gnd 0.58fF
