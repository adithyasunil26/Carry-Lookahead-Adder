magic
tech scmos
timestamp 1618847043
<< metal1 >>
rect -3 1270 97 1273
rect 102 1270 802 1273
rect 3 1263 666 1266
rect 3 1256 6 1263
rect -3 1252 0 1255
rect 241 1212 334 1215
rect 339 1212 533 1215
rect 241 1156 497 1159
rect -3 1153 0 1156
rect -3 1083 0 1086
rect 479 1014 484 1019
rect 494 998 497 1156
rect 530 1148 533 1212
rect 530 1145 549 1148
rect 671 1143 674 1146
rect 897 1137 900 1140
rect 539 1026 542 1036
rect 563 1023 572 1026
rect 970 1001 971 1004
rect 494 995 505 998
rect 563 994 572 997
rect 606 993 618 996
rect 490 989 505 992
rect 566 988 572 991
rect 539 975 542 978
rect 566 966 569 988
rect 495 963 569 966
rect 572 963 576 966
rect 611 939 618 942
rect -3 876 0 879
rect 611 874 614 939
rect 481 871 614 874
rect -3 802 0 805
rect 481 738 484 871
rect 606 762 609 775
rect 568 748 572 751
rect 479 735 484 738
rect 567 742 572 745
rect 630 743 633 746
rect 505 732 509 735
rect 567 734 570 742
rect 563 729 570 734
rect 636 727 643 730
rect 12 718 17 721
rect 636 717 639 727
rect 677 717 680 730
rect 630 714 639 717
rect 606 713 630 714
rect 490 708 507 711
rect 1077 693 1080 696
rect 638 686 643 689
rect 701 685 725 688
rect 487 674 490 682
rect 501 680 507 683
rect 628 680 643 683
rect 487 671 507 674
rect 640 654 643 664
rect 677 661 680 669
rect 627 651 643 654
rect -3 595 0 598
rect 722 551 725 634
rect 480 548 725 551
rect -3 521 0 524
rect 480 457 483 548
rect -3 314 0 317
rect -3 237 0 240
rect -2 30 1 33
rect -2 -8 40 -5
rect 45 -8 569 -5
<< m2contact >>
rect 490 962 495 967
rect 500 732 505 737
rect 633 741 638 746
rect 633 686 638 691
rect 496 680 501 685
<< metal2 >>
rect 481 1199 552 1202
rect 481 1019 484 1199
rect 479 1014 484 1019
rect 481 979 484 987
rect 481 976 504 979
rect 479 735 484 738
rect 12 718 17 721
rect 491 716 494 962
rect 501 737 504 976
rect 491 713 499 716
rect 496 685 499 713
rect 635 691 638 741
<< m123contact >>
rect 97 1270 102 1275
rect 802 1269 807 1274
rect 666 1261 671 1266
rect 334 1212 339 1217
rect 666 1143 671 1148
rect 539 1036 544 1041
rect 742 994 747 999
rect 537 970 542 975
rect 576 963 581 968
rect 549 773 554 778
rect 563 748 568 753
rect 588 651 593 656
rect 40 -9 45 -4
<< metal3 >>
rect 98 1245 101 1270
rect 335 1046 338 1212
rect 667 1148 670 1261
rect 803 1229 806 1269
rect 335 1043 347 1046
rect 344 854 347 1043
rect 407 1043 542 1046
rect 407 1030 410 1043
rect 539 1041 542 1043
rect 667 1041 670 1143
rect 699 1056 702 1164
rect 757 1072 760 1112
rect 757 1069 832 1072
rect 699 1053 775 1056
rect 667 1038 746 1041
rect 743 999 746 1038
rect 772 982 775 1053
rect 829 1034 832 1069
rect 539 966 542 970
rect 539 963 576 966
rect 539 937 542 963
rect 449 934 542 937
rect 344 851 567 854
rect 407 782 553 785
rect 407 749 410 782
rect 550 778 553 782
rect 564 753 567 851
rect 772 806 775 958
rect 876 848 879 912
rect 876 845 939 848
rect 772 803 882 806
rect 879 674 882 803
rect 936 726 939 845
rect 449 653 588 656
rect 41 -4 44 46
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 548 0 1 1105
box -3 -9 349 129
use nor  nor_0
timestamp 1618580541
transform 1 0 505 0 1 1000
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 539 0 1 993
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 572 0 1 999
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1618628987
transform 1 0 621 0 -1 1036
box -3 -9 349 129
use nand  nand_1
timestamp 1618580231
transform 1 0 572 0 -1 740
box 0 -35 34 27
use inv  inv_1
timestamp 1618579805
transform 1 0 606 0 -1 747
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 683
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 643 0 1 691
box 0 -30 34 39
use inv  inv_2
timestamp 1618579805
transform 1 0 677 0 1 684
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1618628987
transform 1 0 728 0 -1 728
box -3 -9 349 129
<< labels >>
rlabel metal1 -3 314 -3 317 3 y3in
rlabel metal1 -3 1153 -3 1156 3 cinin
rlabel metal1 -3 1083 -3 1086 3 x1in
rlabel metal1 -3 876 -3 879 3 y1in
rlabel metal1 -3 802 -3 805 3 x2in
rlabel metal1 -3 595 -3 598 3 y2in
rlabel metal1 -3 521 -3 524 3 x3in
rlabel metal1 -3 237 -3 240 3 x4in
rlabel metal1 -2 30 -2 33 3 y4in
rlabel metal1 -3 1252 -3 1255 3 clk
rlabel metal1 71 1271 71 1271 5 vdd!
rlabel metal1 19 -7 19 -7 1 gnd!
rlabel metal1 900 1137 900 1140 7 z1o
rlabel metal1 971 1001 971 1004 7 z2o
rlabel metal1 1080 693 1080 696 7 z3o
<< end >>
