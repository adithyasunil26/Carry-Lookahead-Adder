* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 vdd a_35_n5# a_30_8# w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=144 ps=60
M1005 a_7_8# a vdd w_n6_2# pfet w=24 l=2
+  ad=144 pd=60 as=0 ps=0
M1006 a_30_n33# a_27_n20# op Gnd nfet w=12 l=2
+  ad=72 pd=36 as=156 ps=50
M1007 op a_11_2# a_7_8# w_n6_2# pfet w=24 l=2
+  ad=312 pd=74 as=0 ps=0
M1008 gnd a_35_n5# a_30_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_7_n33# a gnd Gnd nfet w=12 l=2
+  ad=72 pd=36 as=0 ps=0
M1010 op b a_7_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_30_8# b op w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 m3_n15_10# m2_n15_10# 0.02fF
C1 b m3_n15_10# 0.04fF
C2 w_n6_2# vdd 0.09fF
C3 gnd b 0.13fF
C4 b vdd 0.03fF
C5 m3_n15_10# m1_35_n5# 0.00fF
C6 a a_11_2# 0.04fF
C7 a_35_n5# w_n6_2# 0.06fF
C8 a inv_0/op 0.08fF
C9 m2_35_n5# m3_n15_10# 0.02fF
C10 a_35_n5# b 0.04fF
C11 op m3_n15_10# 0.01fF
C12 a inv_0/w_0_6# 0.08fF
C13 inv_0/w_0_6# inv_0/op 0.04fF
C14 a m3_n15_10# 0.04fF
C15 m3_n15_10# inv_0/op 0.02fF
C16 gnd op 0.04fF
C17 a_35_n5# m1_35_n5# 0.04fF
C18 a_35_n5# a_27_n20# 0.04fF
C19 op vdd 0.03fF
C20 gnd a 0.42fF
C21 a vdd 0.03fF
C22 gnd inv_0/op 0.12fF
C23 inv_0/op vdd 0.15fF
C24 a_35_n5# m2_35_n5# 0.00fF
C25 w_n6_2# inv_1/op 0.08fF
C26 a_35_n5# op 0.06fF
C27 vdd inv_1/w_0_6# 0.06fF
C28 inv_0/w_0_6# vdd 0.06fF
C29 b inv_1/op 0.44fF
C30 a_27_n20# inv_1/op 0.03fF
C31 a_35_n5# m3_n15_10# 0.01fF
C32 w_n6_2# b 0.16fF
C33 op inv_1/op 0.20fF
C34 a_11_2# inv_1/op 0.03fF
C35 a inv_1/op 0.15fF
C36 inv_1/op inv_1/w_0_6# 0.04fF
C37 w_n6_2# op 0.02fF
C38 w_n6_2# a_11_2# 0.08fF
C39 m3_n15_10# inv_1/op 0.25fF
C40 b m2_35_n5# 0.01fF
C41 a w_n6_2# 0.06fF
C42 b op 0.22fF
C43 gnd inv_1/op 0.12fF
C44 a b 0.11fF
C45 inv_0/op m2_n15_10# 0.02fF
C46 vdd inv_1/op 0.15fF
C47 m2_35_n5# m1_35_n5# 0.01fF
C48 op m1_35_n5# 0.07fF
C49 b inv_1/w_0_6# 0.08fF
C50 m3_n15_10# Gnd 0.11fF **FLOATING
C51 m2_35_n5# Gnd 0.08fF **FLOATING
C52 m2_n15_10# Gnd 0.09fF **FLOATING
C53 m1_35_n5# Gnd 0.02fF **FLOATING
C54 a_27_n20# Gnd 0.09fF
C55 op Gnd 0.14fF
C56 a_35_n5# Gnd 0.19fF
C57 a_11_2# Gnd 0.01fF
C58 w_n6_2# Gnd 1.99fF
C59 gnd Gnd 0.39fF
C60 inv_1/op Gnd 0.38fF
C61 b Gnd 1.41fF
C62 inv_1/w_0_6# Gnd 0.58fF
C63 inv_0/op Gnd 0.08fF
C64 vdd Gnd 0.23fF
C65 a Gnd 1.10fF
C66 inv_0/w_0_6# Gnd 0.58fF
