* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 gnd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=5940 pd=3116 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k sumffo_3/xor_0/vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=1080 ps=552
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin sumffo_3/xor_0/vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 sumffo_3/xor_0/vdd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 sumffo_0/xor_0/op cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/op sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k sumffo_3/xor_0/vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 sumffo_0/xor_0/op sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op sumffo_3/xor_0/vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k sumffo_3/xor_0/vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 sumffo_3/xor_0/vdd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 sumffo_2/xor_0/op ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op sumffo_3/xor_0/vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_2/xor_0/op sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 sumffo_1/xor_0/op nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/op sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 sumffo_1/xor_0/op sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 sumffo_3/xor_0/vdd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 sumffo_3/xor_0/op ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/op sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op sumffo_3/xor_0/vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 sumffo_3/xor_0/op sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 gnd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 gnd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd y2in cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 cla_0/l x2in gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_0/l y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 gnd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 gnd y3in cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 cla_0/l x3in gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_0/l y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 gnd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd y2in 1.82fF
C1 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C2 sumffo_3/xor_0/vdd sumffo_2/xor_0/inv_0/op 0.15fF
C3 cla_1/nand_0/a_13_n26# gnd 0.01fF
C4 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C5 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.36fF
C6 x2in ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C7 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C8 cin ffipg_1/k 0.06fF
C9 inv_1/op sumffo_3/xor_0/vdd 0.11fF
C10 sumffo_3/xor_0/vdd sumffo_3/xor_0/a_10_10# 0.93fF
C11 cla_0/nor_1/w_0_0# gnd 0.31fF
C12 x4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C13 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C14 gnd inv_7/w_0_6# 0.15fF
C15 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/xor_0/inv_0/op 0.03fF
C16 cla_0/g0 ffipg_1/k 0.06fF
C17 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C18 cla_2/nand_0/w_0_0# gnd 0.18fF
C19 cin inv_8/w_0_6# 0.06fF
C20 nor_0/a cinbar 0.32fF
C21 sumffo_2/xor_0/inv_0/w_0_6# inv_1/op 0.06fF
C22 gnd nor_4/b 0.25fF
C23 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/op 0.45fF
C24 gnd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C25 gnd sumffo_1/xor_0/a_10_10# 0.93fF
C26 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C27 ffipg_2/k nand_2/b 0.06fF
C28 sumffo_0/xor_0/inv_0/op gnd 0.17fF
C29 gnd inv_5/in 0.49fF
C30 gnd sumffo_1/xor_0/inv_1/op 0.35fF
C31 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C32 gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C33 cla_2/inv_0/in cla_2/p1 0.02fF
C34 inv_2/w_0_6# nor_1/b 0.03fF
C35 cla_2/nor_0/w_0_0# gnd 0.31fF
C36 cla_0/nand_0/w_0_0# cla_0/l 0.06fF
C37 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C38 nor_0/w_0_0# gnd 0.46fF
C39 cla_2/g1 cla_2/inv_0/op 0.35fF
C40 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C41 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C42 gnd nor_2/w_0_0# 0.15fF
C43 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/op 0.52fF
C44 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C45 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C46 inv_5/w_0_6# nor_3/b 0.17fF
C47 x1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C48 gnd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C49 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C50 cla_1/nor_0/w_0_0# gnd 0.31fF
C51 cla_0/g0 cla_0/inv_0/in 0.16fF
C52 cla_0/l y3in 0.13fF
C53 gnd x1in 1.19fF
C54 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C55 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C56 inv_0/in cinbar 0.16fF
C57 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C58 gnd inv_3/in 0.47fF
C59 gnd inv_8/in 0.43fF
C60 cla_2/l cla_0/n 0.32fF
C61 gnd ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C62 inv_1/op ffipg_2/k 0.09fF
C63 inv_9/in cout 0.04fF
C64 nor_2/w_0_0# cla_1/n 0.06fF
C65 inv_1/op nor_1/w_0_0# 0.03fF
C66 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C67 cla_1/p0 gnd 1.12fF
C68 nor_0/w_0_0# inv_0/op 0.10fF
C69 x2in ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C70 inv_7/w_0_6# inv_7/in 0.10fF
C71 x4in ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C72 nand_2/b inv_2/in 0.34fF
C73 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C74 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C75 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C76 cla_2/l inv_7/w_0_6# 0.06fF
C77 cin sumffo_0/xor_0/w_n3_4# 0.06fF
C78 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C79 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C80 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/op 0.02fF
C81 y4in ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C82 nor_3/w_0_0# nor_4/b 0.03fF
C83 gnd cla_1/n 0.52fF
C84 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C85 cin sumffo_1/xor_0/a_10_10# 0.06fF
C86 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# x3in 0.06fF
C87 ffipg_0/pggen_0/nand_0/w_0_0# y1in 0.06fF
C88 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C89 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C90 cla_2/l inv_5/in 0.05fF
C91 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C92 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C93 gnd sumffo_1/xor_0/inv_0/op 0.32fF
C94 inv_0/op gnd 0.27fF
C95 ffipg_0/k nor_0/a 0.05fF
C96 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C97 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C98 y4in ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C99 ffipg_2/k x3in 0.46fF
C100 x2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C101 cin sumffo_0/xor_0/inv_0/op 0.20fF
C102 cin sumffo_1/xor_0/inv_1/op 0.04fF
C103 nor_1/w_0_0# nor_1/b 0.06fF
C104 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C105 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C106 gnd sumffo_2/xor_0/op 0.14fF
C107 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C108 cla_2/g1 y4in 0.13fF
C109 inv_3/w_0_6# nor_2/b 0.03fF
C110 y4in ffipg_3/pggen_0/xor_0/inv_0/op 0.20fF
C111 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.15fF
C112 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C113 nor_0/w_0_0# cin 0.16fF
C114 inv_8/w_0_6# nor_4/a 0.03fF
C115 sumffo_0/xor_0/inv_0/w_0_6# sumffo_3/xor_0/vdd 0.09fF
C116 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.35fF
C117 sumffo_1/xor_0/inv_1/w_0_6# nand_2/b 0.23fF
C118 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C119 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C120 cla_1/inv_0/w_0_6# gnd 0.06fF
C121 sumffo_0/xor_0/w_n3_4# sumffo_3/xor_0/vdd 0.12fF
C122 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C123 nor_0/w_0_0# cla_0/g0 0.06fF
C124 cin sumffo_0/xor_0/a_10_10# 0.12fF
C125 cin sumffo_2/xor_0/w_n3_4# 0.00fF
C126 gnd inv_7/in 0.43fF
C127 gnd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C128 nor_2/w_0_0# inv_4/in 0.11fF
C129 cin inv_8/in 0.13fF
C130 sumffo_0/xor_0/inv_0/op sumffo_3/xor_0/vdd 0.15fF
C131 cla_2/p0 x3in 0.22fF
C132 cla_0/l cla_2/inv_0/in 0.16fF
C133 cla_2/l gnd 0.61fF
C134 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C135 ffipg_1/k nor_0/a 0.06fF
C136 gnd nor_3/w_0_0# 0.14fF
C137 cin gnd 1.19fF
C138 x1in ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C139 cla_2/nor_1/w_0_0# gnd 0.31fF
C140 y3in ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C141 gnd cout 0.25fF
C142 y1in ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C143 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C144 cla_0/g0 cla_1/p0 0.38fF
C145 cla_0/l nand_2/b 0.06fF
C146 inv_6/in nor_4/b 0.04fF
C147 x1in y1in 0.73fF
C148 inv_2/in nor_1/b 0.04fF
C149 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C150 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C151 cla_0/inv_0/op cla_0/l 0.35fF
C152 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C153 nor_4/a inv_9/in 0.02fF
C154 cla_0/g0 gnd 1.23fF
C155 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C156 cla_2/g1 cla_2/nand_0/w_0_0# 0.06fF
C157 nor_4/w_0_0# inv_9/in 0.11fF
C158 cla_2/p1 y4in 0.03fF
C159 gnd inv_4/in 0.33fF
C160 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C161 gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C162 sumffo_3/xor_0/vdd sumffo_0/xor_0/a_10_10# 0.93fF
C163 ffipg_2/k cla_0/n 0.06fF
C164 inv_5/in nor_3/b 0.04fF
C165 ffipg_3/k y4in 0.07fF
C166 y3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C167 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C168 y1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C169 x1in ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C170 nor_1/w_0_0# cla_0/n 0.06fF
C171 sumffo_3/xor_0/vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C172 gnd ffipg_2/pggen_0/nand_0/a_13_n26# 0.01fF
C173 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C174 cla_1/inv_0/op cla_0/n 0.06fF
C175 cin sumffo_1/xor_0/inv_0/op 0.06fF
C176 gnd y1in 1.77fF
C177 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C178 cla_1/nand_0/w_0_0# gnd 0.10fF
C179 gnd inv_2/w_0_6# 0.17fF
C180 y2in ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C181 cin sumffo_2/xor_0/op 0.28fF
C182 sumffo_0/xor_0/inv_1/op ffipg_0/k 0.06fF
C183 gnd sumffo_3/xor_0/vdd 0.75fF
C184 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.32fF
C185 inv_4/in cla_1/n 0.02fF
C186 inv_1/op inv_1/in 0.04fF
C187 inv_0/op cla_0/g0 0.32fF
C188 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C189 y2in ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C190 nor_4/b nor_4/a 0.42fF
C191 ffipg_3/k cla_0/n 0.06fF
C192 nor_4/b nor_4/w_0_0# 0.06fF
C193 x4in y4in 0.73fF
C194 gnd sumffo_3/xor_0/op 0.14fF
C195 sumffo_3/xor_0/vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C196 cla_1/l cla_2/p0 0.02fF
C197 cla_2/inv_0/w_0_6# gnd 0.06fF
C198 gnd cla_2/n 0.60fF
C199 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C200 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C201 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C202 gnd inv_6/in 0.33fF
C203 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.35fF
C204 gnd nor_3/b 0.33fF
C205 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/op 0.02fF
C206 gnd sumffo_1/xor_0/w_n3_4# 0.12fF
C207 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C208 nor_2/b nor_2/w_0_0# 0.06fF
C209 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C210 cla_2/g1 gnd 0.65fF
C211 y3in x3in 0.73fF
C212 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.36fF
C213 y3in ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C214 y1in ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C215 ffipg_0/k cinbar 0.06fF
C216 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C217 cla_1/nor_1/w_0_0# gnd 0.31fF
C218 inv_1/in nor_1/b 0.16fF
C219 sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C220 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C221 inv_3/in nor_2/b 0.04fF
C222 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C223 cla_0/g0 cin 0.08fF
C224 inv_8/in nor_4/a 0.04fF
C225 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C226 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C227 sumffo_3/xor_0/vdd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C228 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C229 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C230 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C231 cla_1/p0 ffipg_2/k 0.06fF
C232 cla_0/inv_0/op nand_2/b 0.09fF
C233 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C234 x2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C235 gnd nor_2/b 0.32fF
C236 cla_1/inv_0/in gnd 0.34fF
C237 gnd nor_4/a 0.40fF
C238 gnd nor_4/w_0_0# 0.15fF
C239 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C240 gnd ffipg_2/k 0.54fF
C241 gnd nor_1/w_0_0# 0.15fF
C242 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/xor_0/inv_0/op 0.03fF
C243 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C244 cla_1/inv_0/op gnd 0.27fF
C245 cin inv_2/w_0_6# 0.06fF
C246 gnd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C247 nor_0/w_0_0# nor_0/a 0.06fF
C248 cin sumffo_3/xor_0/vdd 0.18fF
C249 y2in ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C250 cla_0/g0 y1in 0.13fF
C251 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C252 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.39fF
C253 nor_2/b cla_1/n 0.39fF
C254 sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C255 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C256 cla_2/p1 gnd 1.00fF
C257 cla_0/inv_0/in cla_0/l 0.07fF
C258 cin sumffo_3/xor_0/op 0.16fF
C259 nor_0/a x1in 0.22fF
C260 nor_3/w_0_0# cla_2/n 0.06fF
C261 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/op 0.45fF
C262 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C263 ffipg_1/k x2in 0.46fF
C264 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C265 gnd ffipg_3/k 0.56fF
C266 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C267 cla_2/l nor_3/b 0.10fF
C268 x1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C269 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C270 cla_1/p0 cla_2/p0 0.24fF
C271 nor_3/w_0_0# inv_6/in 0.11fF
C272 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/op 0.52fF
C273 y4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C274 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C275 nor_3/w_0_0# nor_3/b 0.06fF
C276 cla_2/p0 gnd 1.12fF
C277 cin sumffo_1/xor_0/w_n3_4# 0.00fF
C278 cla_1/p0 nor_0/a 0.24fF
C279 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C280 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C281 cla_0/l cla_1/l 0.08fF
C282 y3in ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C283 y1in ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C284 inv_1/in cla_0/n 0.02fF
C285 gnd nor_0/a 0.58fF
C286 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C287 y2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C288 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C289 gnd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C290 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/op 0.02fF
C291 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C292 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C293 gnd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C294 cla_0/l cla_0/n 0.25fF
C295 nor_0/w_0_0# inv_0/in 0.11fF
C296 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C297 gnd inv_2/in 0.47fF
C298 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C299 sumffo_2/xor_0/inv_1/w_0_6# ffipg_2/k 0.23fF
C300 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C301 gnd x4in 1.24fF
C302 cla_0/l y2in 0.13fF
C303 ffipg_3/pggen_0/nand_0/w_0_0# y4in 0.06fF
C304 sumffo_2/xor_0/inv_0/w_0_6# sumffo_3/xor_0/vdd 0.09fF
C305 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/op 0.06fF
C306 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C307 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C308 sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_0/op 0.15fF
C309 inv_1/op sumffo_2/xor_0/inv_0/op 0.27fF
C310 ffipg_1/k nand_2/b 0.15fF
C311 cla_0/l inv_7/w_0_6# 0.06fF
C312 gnd sumffo_1/xor_0/op 0.14fF
C313 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C314 nor_4/w_0_0# cout 0.03fF
C315 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C316 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/op 0.06fF
C317 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C318 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C319 nand_2/b inv_3/w_0_6# 0.06fF
C320 gnd inv_0/in 0.30fF
C321 inv_6/in cla_2/n 0.02fF
C322 cla_0/nand_0/a_13_n26# gnd 0.00fF
C323 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.36fF
C324 nor_2/b inv_4/in 0.16fF
C325 cla_2/n nor_3/b 0.41fF
C326 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/op 0.45fF
C327 gnd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C328 cla_2/l cla_2/p1 0.02fF
C329 cla_2/g1 cla_2/n 0.13fF
C330 cla_0/nand_0/w_0_0# gnd 0.10fF
C331 y2in x2in 0.73fF
C332 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C333 inv_6/in nor_3/b 0.16fF
C334 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C335 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C336 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C337 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C338 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/op 0.06fF
C339 gnd sumffo_0/xor_0/op 0.14fF
C340 cla_2/l cla_2/p0 0.16fF
C341 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C342 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C343 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C344 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C345 sumffo_3/xor_0/vdd ffipg_2/k 0.10fF
C346 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C347 gnd y3in 1.82fF
C348 inv_0/op inv_0/in 0.04fF
C349 inv_7/op inv_8/w_0_6# 0.06fF
C350 cla_2/nand_0/a_13_n26# gnd 0.01fF
C351 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C352 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C353 inv_4/op nor_2/w_0_0# 0.03fF
C354 gnd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C355 gnd inv_1/in 0.33fF
C356 x2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C357 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C358 cla_0/l cla_1/p0 0.09fF
C359 cla_1/l nand_2/b 0.31fF
C360 cin inv_2/in 0.13fF
C361 cla_0/l gnd 3.30fF
C362 cla_0/g0 nor_0/a 0.57fF
C363 nor_0/w_0_0# cinbar 0.06fF
C364 x2in ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C365 nand_2/b cla_0/n 0.06fF
C366 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C367 sumffo_3/xor_0/vdd ffipg_3/k 0.10fF
C368 cla_0/nor_0/w_0_0# gnd 0.31fF
C369 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C370 gnd inv_4/op 0.47fF
C371 nor_0/a y1in 0.03fF
C372 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C373 cin sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C374 cin sumffo_1/xor_0/op 0.27fF
C375 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C376 x3in ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C377 y1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C378 cla_0/l cla_1/n 0.13fF
C379 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C380 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C381 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C382 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C383 cin inv_0/in 0.07fF
C384 inv_2/w_0_6# inv_2/in 0.10fF
C385 gnd cinbar 0.16fF
C386 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C387 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C388 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C389 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C390 y4in ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C391 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C392 cla_1/p0 x2in 0.22fF
C393 cla_2/g1 cla_2/p1 0.00fF
C394 cin sumffo_1/xor_0/a_38_n43# 0.01fF
C395 gnd x2in 1.24fF
C396 nor_4/a nor_4/w_0_0# 0.07fF
C397 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C398 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C399 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C400 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C401 ffipg_2/pggen_0/nand_0/w_0_0# y3in 0.06fF
C402 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C403 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C404 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C405 inv_7/op inv_7/w_0_6# 0.03fF
C406 nor_0/w_0_0# nand_2/b 0.04fF
C407 y2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C408 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C409 sumffo_0/xor_0/inv_1/w_0_6# sumffo_3/xor_0/vdd 0.06fF
C410 sumffo_3/xor_0/inv_0/w_0_6# inv_4/op 0.06fF
C411 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C412 cla_0/l inv_7/in 0.13fF
C413 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C414 cla_0/n inv_5/w_0_6# 0.06fF
C415 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C416 cin sumffo_0/xor_0/inv_1/op 0.22fF
C417 cla_2/inv_0/in gnd 0.34fF
C418 cla_2/l cla_0/l 0.37fF
C419 x4in ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C420 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C421 nand_2/b inv_3/in 0.13fF
C422 cla_0/l cin 0.33fF
C423 cla_2/inv_0/op cla_2/nand_0/w_0_0# 0.06fF
C424 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C425 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/op 0.45fF
C426 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C427 cla_1/inv_0/in cla_2/p0 0.02fF
C428 cla_0/inv_0/w_0_6# gnd 0.06fF
C429 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.11fF
C430 cla_2/p0 ffipg_2/k 0.05fF
C431 nor_1/b cla_0/n 0.36fF
C432 gnd nand_2/b 1.92fF
C433 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/op 0.02fF
C434 gnd ffipg_1/pggen_0/nand_0/a_13_n26# 0.01fF
C435 ffipg_1/k y2in 0.07fF
C436 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op 0.52fF
C437 cla_0/inv_0/op gnd 0.27fF
C438 cla_1/l inv_3/w_0_6# 0.06fF
C439 cla_0/g0 cla_0/l 0.14fF
C440 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C441 x3in ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C442 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C443 inv_3/w_0_6# cla_0/n 0.16fF
C444 cla_2/p1 ffipg_3/k 0.05fF
C445 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_1/op 0.08fF
C446 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C447 gnd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C448 ffipg_0/k x1in 0.46fF
C449 inv_5/w_0_6# inv_5/in 0.10fF
C450 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C451 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C452 cla_2/p0 cla_2/p1 0.24fF
C453 cin sumffo_2/xor_0/a_38_n43# 0.01fF
C454 inv_4/op inv_4/in 0.04fF
C455 sumffo_0/xor_0/inv_1/op sumffo_3/xor_0/vdd 0.15fF
C456 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C457 cla_0/l inv_2/w_0_6# 0.06fF
C458 cla_2/p0 ffipg_3/k 0.06fF
C459 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C460 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C461 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C462 inv_7/op gnd 0.27fF
C463 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C464 cin sumffo_2/xor_0/a_10_10# 0.04fF
C465 gnd ffipg_0/k 0.57fF
C466 gnd sumffo_2/xor_0/inv_0/op 0.17fF
C467 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C468 cla_2/p1 x4in 0.22fF
C469 y2in ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C470 cin sumffo_2/xor_0/inv_1/op 0.04fF
C471 inv_1/op gnd 0.47fF
C472 sumffo_3/xor_0/vdd inv_4/op 0.11fF
C473 ffipg_3/k x4in 0.46fF
C474 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.15fF
C475 cla_2/inv_0/op gnd 0.27fF
C476 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C477 cla_1/l cla_0/n 0.07fF
C478 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C479 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C480 gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C481 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C482 gnd inv_5/w_0_6# 0.42fF
C483 cla_0/l cla_2/g1 0.26fF
C484 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C485 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C486 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C487 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C488 cin sumffo_3/xor_0/inv_1/op 0.04fF
C489 y1in ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C490 sumffo_3/xor_0/vdd sumffo_2/xor_0/a_10_10# 0.93fF
C491 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C492 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C493 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op 0.06fF
C494 ffipg_2/k y3in 0.07fF
C495 cla_1/p0 ffipg_1/k 0.05fF
C496 cin nand_2/b 0.04fF
C497 gnd ffipg_0/pggen_0/nand_0/a_13_n26# 0.01fF
C498 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C499 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C500 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C501 gnd ffipg_1/k 0.76fF
C502 sumffo_3/xor_0/vdd sumffo_2/xor_0/inv_1/op 0.15fF
C503 gnd x3in 1.24fF
C504 gnd nor_1/b 0.35fF
C505 inv_3/w_0_6# inv_3/in 0.10fF
C506 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.39fF
C507 nor_1/w_0_0# inv_1/in 0.11fF
C508 inv_8/w_0_6# inv_8/in 0.10fF
C509 nor_4/b inv_9/in 0.16fF
C510 cla_0/l cla_1/inv_0/in 0.23fF
C511 inv_7/op inv_7/in 0.04fF
C512 cla_0/g0 nand_2/b 0.13fF
C513 inv_0/in nor_0/a 0.02fF
C514 cla_0/l ffipg_2/k 0.10fF
C515 gnd inv_3/w_0_6# 0.17fF
C516 gnd inv_8/w_0_6# 0.15fF
C517 cla_0/l cla_1/inv_0/op 0.35fF
C518 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C519 y2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C520 cla_0/n inv_5/in 0.13fF
C521 inv_7/op cin 0.31fF
C522 sumffo_3/xor_0/vdd sumffo_3/xor_0/inv_1/op 0.15fF
C523 ffipg_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C524 nand_2/b inv_2/w_0_6# 0.03fF
C525 cin ffipg_0/k 0.19fF
C526 cin sumffo_2/xor_0/inv_0/op 0.06fF
C527 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C528 cla_0/inv_0/in cla_1/p0 0.02fF
C529 cin sumffo_3/xor_0/a_38_n43# 0.01fF
C530 cla_2/p0 y3in 0.03fF
C531 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C532 gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C533 cla_0/l cla_2/p1 0.30fF
C534 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C535 cla_0/inv_0/in gnd 0.34fF
C536 gnd y4in 1.76fF
C537 cla_0/l ffipg_3/k 0.10fF
C538 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/op 0.52fF
C539 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C540 cin sumffo_3/xor_0/a_10_10# 0.04fF
C541 x3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C542 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C543 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C544 ffipg_0/pggen_0/nand_0/w_0_0# x1in 0.06fF
C545 cla_0/l cla_2/p0 0.44fF
C546 cla_1/p0 cla_1/l 0.16fF
C547 cla_2/l inv_5/w_0_6# 0.08fF
C548 cla_2/g1 cla_2/inv_0/in 0.04fF
C549 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C550 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C551 inv_4/op ffipg_3/k 0.09fF
C552 cla_1/l gnd 0.40fF
C553 ffipg_0/k y1in 0.07fF
C554 cla_0/l nor_0/a 0.16fF
C555 gnd inv_9/in 0.33fF
C556 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C557 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C558 y4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C559 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C560 cla_1/p0 y2in 0.03fF
C561 gnd cla_0/n 1.18fF
C562 ffipg_2/pggen_0/nand_0/w_0_0# x3in 0.06fF
C563 gnd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C564 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C565 ffipg_0/k sumffo_3/xor_0/vdd 0.11fF
C566 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C567 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C568 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C569 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C570 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C571 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C572 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C573 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C574 y4in Gnd 2.72fF
C575 x4in Gnd 2.80fF
C576 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C577 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C578 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C579 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C580 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C581 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C582 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C583 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C584 y3in Gnd 2.72fF
C585 x3in Gnd 2.80fF
C586 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C587 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C588 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C589 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C590 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C591 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C592 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C593 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C594 y2in Gnd 2.72fF
C595 x2in Gnd 2.80fF
C596 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C597 cout Gnd 0.19fF
C598 inv_9/in Gnd 0.23fF
C599 nor_4/w_0_0# Gnd 1.81fF
C600 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C601 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C602 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C603 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C604 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C605 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C606 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C607 y1in Gnd 2.72fF
C608 x1in Gnd 2.80fF
C609 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C610 nor_4/a Gnd 0.59fF
C611 inv_8/in Gnd 0.22fF
C612 inv_8/w_0_6# Gnd 1.40fF
C613 inv_7/in Gnd 0.22fF
C614 inv_7/w_0_6# Gnd 1.40fF
C615 nor_4/b Gnd 0.32fF
C616 nor_3/b Gnd 0.77fF
C617 inv_5/in Gnd 0.22fF
C618 inv_5/w_0_6# Gnd 1.40fF
C619 cla_2/n Gnd 0.36fF
C620 inv_6/in Gnd 0.23fF
C621 nor_3/w_0_0# Gnd 1.81fF
C622 cla_1/n Gnd 0.36fF
C623 inv_4/in Gnd 0.23fF
C624 nor_2/w_0_0# Gnd 1.81fF
C625 cla_0/n Gnd 1.34fF
C626 nor_2/b Gnd 0.82fF
C627 inv_3/in Gnd 0.22fF
C628 inv_3/w_0_6# Gnd 1.40fF
C629 cinbar Gnd 1.21fF
C630 nor_0/a Gnd 2.07fF
C631 nor_1/b Gnd 1.05fF
C632 inv_2/in Gnd 0.22fF
C633 inv_2/w_0_6# Gnd 1.40fF
C634 inv_1/in Gnd 0.23fF
C635 nor_1/w_0_0# Gnd 1.81fF
C636 inv_0/in Gnd 0.23fF
C637 sumffo_3/xor_0/op Gnd 0.06fF
C638 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C639 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C640 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C641 ffipg_3/k Gnd 2.89fF
C642 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C643 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C644 inv_4/op Gnd 1.37fF
C645 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C646 sumffo_1/xor_0/op Gnd 0.06fF
C647 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C648 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C649 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C650 nand_2/b Gnd 2.33fF
C651 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C652 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C653 ffipg_1/k Gnd 2.78fF
C654 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C655 sumffo_2/xor_0/op Gnd 0.06fF
C656 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C657 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C658 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C659 ffipg_2/k Gnd 2.89fF
C660 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C661 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C662 inv_1/op Gnd 1.30fF
C663 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C664 sumffo_0/xor_0/op Gnd 0.06fF
C665 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C666 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C667 gnd Gnd 29.42fF
C668 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C669 sumffo_3/xor_0/vdd Gnd 1.76fF
C670 cin Gnd 7.80fF
C671 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C672 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C673 ffipg_0/k Gnd 1.49fF
C674 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C675 cla_2/p1 Gnd 1.09fF
C676 cla_2/nor_1/w_0_0# Gnd 1.23fF
C677 cla_2/nor_0/w_0_0# Gnd 1.23fF
C678 cla_2/inv_0/in Gnd 0.27fF
C679 cla_2/inv_0/w_0_6# Gnd 0.58fF
C680 cla_2/g1 Gnd 0.59fF
C681 cla_2/inv_0/op Gnd 0.26fF
C682 cla_2/nand_0/w_0_0# Gnd 0.82fF
C683 cla_2/p0 Gnd 0.38fF
C684 cla_1/nor_1/w_0_0# Gnd 1.23fF
C685 cla_1/l Gnd 0.30fF
C686 cla_1/nor_0/w_0_0# Gnd 1.23fF
C687 cla_1/inv_0/in Gnd 0.27fF
C688 cla_1/inv_0/w_0_6# Gnd 0.58fF
C689 cla_1/inv_0/op Gnd 0.26fF
C690 cla_1/nand_0/w_0_0# Gnd 0.82fF
C691 inv_7/op Gnd 0.26fF
C692 cla_1/p0 Gnd 2.28fF
C693 cla_0/nor_1/w_0_0# Gnd 1.23fF
C694 cla_0/l Gnd 3.41fF
C695 cla_0/nor_0/w_0_0# Gnd 1.23fF
C696 cla_0/inv_0/in Gnd 0.27fF
C697 cla_0/inv_0/w_0_6# Gnd 0.58fF
C698 cla_0/inv_0/op Gnd 0.26fF
C699 cla_0/nand_0/w_0_0# Gnd 0.82fF
C700 cla_2/l Gnd 0.25fF
C701 cla_0/g0 Gnd 1.40fF
C702 inv_0/op Gnd 0.23fF
C703 nor_0/w_0_0# Gnd 2.63fF
