magic
tech scmos
timestamp 1619548844
<< metal1 >>
rect 324 1511 391 1514
rect 396 1511 523 1514
rect 528 1511 627 1514
rect 632 1511 727 1514
rect 324 1487 561 1490
rect 558 1434 561 1487
rect 601 1460 615 1463
rect 601 1436 604 1460
rect 731 1441 733 1444
rect 324 1431 510 1434
rect 472 1309 475 1405
rect 507 1363 510 1431
rect 558 1431 599 1434
rect 558 1425 561 1431
rect 531 1406 615 1409
rect 507 1360 516 1363
rect 247 1291 249 1294
rect 513 1291 516 1360
rect 553 1329 558 1332
rect 555 1319 558 1329
rect 611 1316 617 1319
rect 652 1302 654 1305
rect 513 1288 519 1291
rect 611 1286 612 1289
rect 617 1286 642 1289
rect 472 1282 501 1285
rect 506 1282 519 1285
rect 550 1263 553 1274
rect 472 1256 494 1259
rect 499 1256 565 1259
rect 574 1257 577 1271
rect 758 1267 760 1270
rect 611 1257 620 1260
rect 248 1237 250 1240
rect 634 1232 642 1235
rect 634 1171 637 1232
rect 472 1168 637 1171
rect 472 1068 475 1168
rect 613 1097 616 1108
rect 576 1081 579 1084
rect 572 1075 579 1078
rect 637 1076 640 1079
rect 508 1065 509 1068
rect 572 1065 575 1075
rect 568 1062 575 1065
rect 247 1050 249 1053
rect 641 1050 648 1053
rect 637 1047 644 1050
rect 611 1046 637 1047
rect 472 1041 487 1044
rect 492 1041 507 1044
rect 682 1040 685 1053
rect 469 1007 472 1015
rect 501 1013 507 1016
rect 625 1008 628 1013
rect 644 1009 648 1012
rect 706 1008 714 1011
rect 469 1004 476 1007
rect 481 1004 507 1007
rect 630 1003 648 1006
rect 248 996 250 999
rect 706 993 726 996
rect 706 992 709 993
rect 627 984 648 987
rect 682 984 685 992
rect 830 973 832 976
rect 694 954 714 957
rect 694 940 697 954
rect 472 937 548 940
rect 552 937 697 940
rect 472 849 475 937
rect 609 878 612 889
rect 568 862 575 865
rect 570 856 575 859
rect 632 857 635 860
rect 494 846 507 849
rect 570 846 573 856
rect 568 843 573 846
rect 247 831 249 834
rect 641 831 647 834
rect 632 828 644 831
rect 609 827 633 828
rect 472 822 499 825
rect 504 822 507 825
rect 681 821 684 834
rect 469 788 472 796
rect 480 794 507 797
rect 469 785 479 788
rect 484 785 507 788
rect 625 787 628 794
rect 641 790 647 793
rect 705 789 711 792
rect 625 784 647 787
rect 248 777 250 780
rect 705 774 723 777
rect 705 773 708 774
rect 627 765 647 768
rect 681 765 684 773
rect 827 754 829 757
rect 695 735 711 738
rect 695 716 698 735
rect 472 713 698 716
rect 472 626 475 713
rect 631 667 655 670
rect 607 655 610 666
rect 631 650 634 667
rect 685 657 688 670
rect 715 657 718 671
rect 752 658 755 671
rect 709 654 718 657
rect 648 643 651 646
rect 568 639 573 642
rect 645 639 651 640
rect 567 633 573 636
rect 648 637 651 639
rect 709 638 718 641
rect 567 623 570 633
rect 565 620 570 623
rect 247 608 249 611
rect 709 609 718 612
rect 752 609 755 610
rect 685 608 688 609
rect 631 605 638 608
rect 607 604 631 605
rect 472 599 504 602
rect 672 595 675 608
rect 696 592 705 595
rect 739 582 742 595
rect 469 565 472 573
rect 484 571 504 574
rect 469 562 504 565
rect 622 561 625 571
rect 782 569 787 572
rect 634 564 638 567
rect 696 563 702 566
rect 622 558 638 561
rect 248 554 250 557
rect 699 554 702 563
rect 699 551 705 554
rect 782 553 785 569
rect 763 550 785 553
rect 607 519 610 542
rect 621 539 638 542
rect 672 539 675 547
rect 693 529 696 547
rect 693 526 705 529
rect 739 526 742 534
rect 268 516 297 519
rect 302 516 799 519
<< m2contact >>
rect 472 1405 477 1410
rect 557 1420 562 1425
rect 526 1406 531 1411
rect 647 1301 652 1306
rect 612 1285 617 1290
rect 501 1280 506 1285
rect 575 1279 580 1284
rect 494 1255 499 1260
rect 565 1256 570 1261
rect 620 1257 625 1262
rect 571 1081 576 1086
rect 640 1076 645 1081
rect 503 1065 508 1070
rect 487 1039 492 1044
rect 496 1013 501 1018
rect 639 1009 644 1014
rect 476 1003 481 1008
rect 625 1003 630 1008
rect 563 862 568 867
rect 489 846 494 851
rect 635 855 640 860
rect 499 820 504 825
rect 475 794 480 799
rect 479 783 484 788
rect 636 790 641 795
rect 607 650 612 655
rect 563 639 568 644
rect 629 634 634 639
rect 499 623 504 628
rect 479 571 484 576
rect 629 564 634 569
rect 605 542 610 547
<< metal2 >>
rect 477 1407 526 1410
rect 477 799 480 1003
rect 489 851 492 1039
rect 496 1018 499 1255
rect 503 1070 506 1280
rect 519 1111 522 1332
rect 558 1084 561 1420
rect 648 1306 651 1364
rect 622 1302 647 1305
rect 575 1261 578 1279
rect 570 1258 578 1261
rect 612 1117 615 1285
rect 622 1262 625 1302
rect 601 1114 615 1117
rect 558 1081 571 1084
rect 519 892 522 970
rect 601 947 604 1114
rect 640 1014 643 1076
rect 563 944 604 947
rect 563 867 566 944
rect 627 921 630 1003
rect 579 918 630 921
rect 481 576 484 783
rect 501 628 504 820
rect 520 747 523 751
rect 517 744 523 747
rect 517 669 520 744
rect 579 680 582 918
rect 636 795 639 855
rect 563 677 582 680
rect 563 644 566 677
rect 609 655 612 765
rect 607 547 610 650
rect 629 569 632 634
<< m123contact >>
rect 391 1511 396 1516
rect 523 1511 528 1516
rect 627 1511 632 1516
rect 599 1431 604 1436
rect 522 1329 527 1334
rect 647 1364 652 1369
rect 617 1315 622 1320
rect 599 1255 604 1260
rect 546 1062 551 1067
rect 613 1092 618 1097
rect 701 1037 706 1042
rect 611 982 616 987
rect 609 873 614 878
rect 700 818 705 823
rect 609 765 614 770
rect 559 620 564 625
rect 643 643 648 648
rect 713 644 718 649
rect 773 639 778 644
rect 643 634 648 639
rect 700 543 705 548
rect 297 514 302 519
<< metal3 >>
rect 392 1323 395 1511
rect 524 1334 527 1511
rect 628 1432 631 1511
rect 601 1357 604 1431
rect 647 1369 650 1423
rect 601 1354 737 1357
rect 622 1316 634 1319
rect 298 1227 307 1230
rect 304 989 307 1227
rect 298 986 307 989
rect 283 768 295 771
rect 304 770 307 986
rect 283 594 286 768
rect 298 767 307 770
rect 441 606 444 1294
rect 631 1258 634 1316
rect 631 1255 654 1258
rect 600 1136 603 1255
rect 600 1133 616 1136
rect 613 1097 616 1133
rect 734 1101 737 1354
rect 734 1098 809 1101
rect 548 1019 551 1062
rect 548 1016 600 1019
rect 597 686 600 1016
rect 613 987 616 1092
rect 706 1039 726 1042
rect 611 878 614 982
rect 610 770 613 873
rect 705 819 723 822
rect 806 697 809 1098
rect 713 694 809 697
rect 596 683 646 686
rect 643 648 646 683
rect 713 649 716 694
rect 643 623 646 634
rect 564 620 646 623
rect 778 603 781 642
rect 702 600 781 603
rect 702 548 705 600
rect 297 519 300 544
use sumffo  sumffo_0
timestamp 1619451829
transform 1 0 618 0 -1 1503
box -3 24 113 129
use ffipg  ffipg_0
timestamp 1619450786
transform 1 0 2 0 1 1139
box 247 76 470 193
use nor  nor_0
timestamp 1618580541
transform 1 0 519 0 1 1293
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 553 0 1 1286
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 577 0 1 1292
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1619451829
transform 1 0 645 0 -1 1329
box -3 24 113 129
use ffipg  ffipg_1
timestamp 1619450786
transform 1 0 2 0 1 898
box 247 76 470 193
use nand  nand_1
timestamp 1618580231
transform 1 0 579 0 -1 1073
box 0 -35 34 27
use inv  inv_2
timestamp 1618579805
transform 1 0 613 0 -1 1080
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 1016
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 648 0 1 1014
box 0 -30 34 39
use inv  inv_1
timestamp 1618579805
transform 1 0 682 0 1 1007
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1619451829
transform 1 0 717 0 1 914
box -3 24 113 129
use ffipg  ffipg_2
timestamp 1619450786
transform 1 0 2 0 1 679
box 247 76 470 193
use nand  nand_2
timestamp 1618580231
transform 1 0 575 0 -1 854
box 0 -35 34 27
use inv  inv_3
timestamp 1618579805
transform 1 0 609 0 -1 861
box 0 -15 24 33
use cla  cla_1
timestamp 1618627066
transform 1 0 516 0 1 797
box -9 -46 112 95
use nor  nor_2
timestamp 1618580541
transform 1 0 647 0 1 795
box 0 -30 34 39
use inv  inv_4
timestamp 1618579805
transform 1 0 681 0 1 788
box 0 -15 24 33
use sumffo  sumffo_3
timestamp 1619451829
transform 1 0 714 0 1 695
box -3 24 113 129
use ffipg  ffipg_3
timestamp 1619450786
transform 1 0 2 0 1 456
box 247 76 470 193
use nand  nand_3
timestamp 1618580231
transform 1 0 573 0 -1 631
box 0 -35 34 27
use inv  inv_5
timestamp 1618579805
transform 1 0 607 0 -1 638
box 0 -15 24 33
use nand  nand_4
timestamp 1618580231
transform 1 0 651 0 -1 635
box 0 -35 34 27
use inv  inv_7
timestamp 1618579805
transform 1 0 685 0 -1 642
box 0 -15 24 33
use nand  nand_5
timestamp 1618580231
transform 1 0 718 0 -1 636
box 0 -35 34 27
use inv  inv_8
timestamp 1618579805
transform 1 0 752 0 -1 643
box 0 -15 24 33
use cla  cla_2
timestamp 1618627066
transform 1 0 513 0 1 574
box -9 -46 112 95
use nor  nor_3
timestamp 1618580541
transform 1 0 638 0 1 569
box 0 -30 34 39
use inv  inv_6
timestamp 1618579805
transform 1 0 672 0 1 562
box 0 -15 24 33
use nor  nor_4
timestamp 1618580541
transform 1 0 705 0 1 556
box 0 -30 34 39
use inv  inv_9
timestamp 1618579805
transform 1 0 739 0 1 549
box 0 -15 24 33
<< labels >>
rlabel metal1 247 831 247 834 3 x3in
rlabel metal1 248 777 248 780 3 y3in
rlabel metal1 247 608 247 611 3 x4in
rlabel metal1 248 554 248 557 3 y4in
rlabel metal1 787 569 787 572 1 cout
rlabel metal1 311 517 311 517 1 gnd!
rlabel metal1 247 1050 247 1053 3 x2in
rlabel metal1 248 996 248 999 3 y2in
rlabel metal1 247 1291 247 1294 3 x1in
rlabel metal1 248 1237 248 1240 3 y1in
rlabel metal1 506 1512 506 1512 5 vdd!
rlabel metal1 324 1487 324 1490 1 cin
rlabel metal1 324 1431 324 1434 1 cinbar
rlabel metal1 832 973 832 976 7 s3
rlabel metal1 760 1267 760 1270 1 s2
rlabel metal1 733 1441 733 1444 1 s1
rlabel metal1 829 754 829 757 7 s4
<< end >>
