* SPICE3 file created from sumffo.ext - technology: scmos

.option scale=0.09u

M1000 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=720 ps=428
M1001 vdd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=1440 pd=796 as=96 ps=40
M1002 ffo_0/nand_3/b ffo_0/nand_1/a vdd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 ffo_0/nand_1/a ffo_0/inv_0/op vdd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 ffo_0/nand_3/a ffo_0/d vdd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 ffo_0/nand_1/b ffo_0/nand_3/a vdd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 ffo_0/nand_6/a ffo_0/nand_3/b vdd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 ffo_0/nand_7/a clk vdd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1025 vdd s sbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1026 sbar ffo_0/nand_6/a vdd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 sbar s ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1028 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1029 vdd sbar s ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1030 s ffo_0/nand_7/a vdd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 s sbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1032 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1033 ffo_0/inv_0/op ffo_0/d vdd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1034 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1035 ffo_0/nand_0/b clk vdd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1036 xor_0/inv_0/op k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1037 xor_0/inv_0/op k vdd xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 xor_0/inv_1/op c gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1039 xor_0/inv_1/op c vdd xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1040 vdd c xor_0/a_10_10# xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1041 ffo_0/d c xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1042 gnd xor_0/inv_1/op xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1043 xor_0/a_10_10# xor_0/inv_1/op ffo_0/d xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1044 xor_0/a_10_n43# k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 xor_0/a_38_n43# xor_0/inv_0/op ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 xor_0/a_10_10# k vdd xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 ffo_0/d xor_0/inv_0/op xor_0/a_10_10# xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ffo_0/d xor_0/inv_0/op 0.06fF
C1 xor_0/inv_0/w_0_6# k 0.06fF
C2 clk vdd 1.49fF
C3 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C4 xor_0/inv_0/op vdd 0.15fF
C5 ffo_0/nand_5/w_0_0# clk 0.06fF
C6 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C7 xor_0/inv_0/w_0_6# vdd 0.09fF
C8 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C9 ffo_0/nand_7/w_0_0# s 0.04fF
C10 ffo_0/nand_0/b clk 0.04fF
C11 vdd xor_0/inv_1/w_0_6# 0.06fF
C12 ffo_0/nand_1/b vdd 0.31fF
C13 xor_0/inv_1/op xor_0/inv_0/op 0.08fF
C14 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C15 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C16 ffo_0/nand_3/a gnd 0.03fF
C17 xor_0/inv_0/w_0_6# xor_0/inv_0/op 0.03fF
C18 ffo_0/nand_7/a s 0.00fF
C19 xor_0/inv_1/op xor_0/inv_1/w_0_6# 0.03fF
C20 ffo_0/nand_3/b gnd 0.35fF
C21 xor_0/w_n3_4# xor_0/a_10_10# 0.16fF
C22 ffo_0/d xor_0/a_10_10# 0.45fF
C23 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C24 clk ffo_0/nand_1/b 0.45fF
C25 ffo_0/nand_4/w_0_0# vdd 0.10fF
C26 ffo_0/nand_3/w_0_0# ffo_0/nand_3/a 0.06fF
C27 vdd xor_0/a_10_10# 0.93fF
C28 ffo_0/nand_3/w_0_0# ffo_0/nand_3/b 0.06fF
C29 ffo_0/nand_7/a gnd 0.03fF
C30 ffo_0/nand_3/a vdd 0.30fF
C31 c gnd 0.11fF
C32 vdd ffo_0/nand_7/w_0_0# 0.10fF
C33 ffo_0/nand_3/b vdd 0.39fF
C34 ffo_0/nand_4/w_0_0# clk 0.06fF
C35 ffo_0/nand_1/w_0_0# ffo_0/nand_1/a 0.06fF
C36 ffo_0/nand_0/b ffo_0/nand_3/a 0.13fF
C37 k c 0.09fF
C38 xor_0/w_n3_4# c 0.06fF
C39 sbar ffo_0/nand_7/w_0_0# 0.06fF
C40 ffo_0/nand_6/w_0_0# s 0.06fF
C41 vdd ffo_0/nand_7/a 0.30fF
C42 c vdd 0.10fF
C43 ffo_0/nand_6/w_0_0# ffo_0/nand_6/a 0.06fF
C44 ffo_0/nand_5/w_0_0# ffo_0/nand_7/a 0.04fF
C45 ffo_0/nand_3/b clk 0.33fF
C46 ffo_0/nand_1/w_0_0# vdd 0.10fF
C47 vdd ffo_0/inv_1/w_0_6# 0.06fF
C48 sbar ffo_0/nand_7/a 0.31fF
C49 ffo_0/nand_6/a s 0.31fF
C50 ffo_0/inv_0/op gnd 0.10fF
C51 xor_0/inv_1/op c 0.22fF
C52 xor_0/inv_0/op c 0.20fF
C53 ffo_0/nand_3/b ffo_0/nand_1/b 0.32fF
C54 ffo_0/nand_0/b ffo_0/inv_1/w_0_6# 0.03fF
C55 s gnd 0.52fF
C56 ffo_0/d ffo_0/inv_0/op 0.04fF
C57 clk ffo_0/inv_1/w_0_6# 0.06fF
C58 ffo_0/nand_6/a gnd 0.03fF
C59 c xor_0/inv_1/w_0_6# 0.23fF
C60 ffo_0/nand_6/w_0_0# vdd 0.10fF
C61 ffo_0/nand_1/b ffo_0/nand_7/a 0.13fF
C62 ffo_0/inv_0/op vdd 0.17fF
C63 ffo_0/inv_0/op ffo_0/nand_0/w_0_0# 0.06fF
C64 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C65 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C66 ffo_0/nand_0/b ffo_0/inv_0/op 0.32fF
C67 ffo_0/nand_1/a gnd 0.03fF
C68 vdd s 0.28fF
C69 ffo_0/inv_0/op ffo_0/inv_0/w_0_6# 0.03fF
C70 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C71 ffo_0/nand_6/w_0_0# sbar 0.04fF
C72 ffo_0/nand_6/a vdd 0.30fF
C73 k gnd 0.22fF
C74 ffo_0/nand_2/w_0_0# ffo_0/d 0.06fF
C75 c xor_0/a_10_10# 0.12fF
C76 ffo_0/d gnd 0.37fF
C77 ffo_0/nand_2/w_0_0# vdd 0.10fF
C78 vdd gnd 0.28fF
C79 ffo_0/nand_7/w_0_0# ffo_0/nand_7/a 0.06fF
C80 sbar s 0.32fF
C81 ffo_0/nand_6/a sbar 0.00fF
C82 ffo_0/nand_1/a vdd 0.30fF
C83 ffo_0/nand_1/a ffo_0/nand_0/w_0_0# 0.04fF
C84 clk ffo_0/nand_6/a 0.13fF
C85 xor_0/w_n3_4# k 0.06fF
C86 ffo_0/d xor_0/w_n3_4# 0.02fF
C87 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C88 ffo_0/nand_3/w_0_0# vdd 0.11fF
C89 ffo_0/nand_0/b gnd 0.38fF
C90 k vdd 0.11fF
C91 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C92 xor_0/w_n3_4# vdd 0.12fF
C93 ffo_0/nand_0/b ffo_0/nand_1/a 0.13fF
C94 ffo_0/d vdd 0.04fF
C95 xor_0/inv_1/op gnd 0.20fF
C96 sbar gnd 0.34fF
C97 clk gnd 0.17fF
C98 ffo_0/nand_0/w_0_0# vdd 0.10fF
C99 xor_0/inv_0/op gnd 0.17fF
C100 ffo_0/nand_5/w_0_0# vdd 0.10fF
C101 ffo_0/d ffo_0/nand_0/b 0.40fF
C102 xor_0/inv_1/op k 0.06fF
C103 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C104 xor_0/inv_1/op xor_0/w_n3_4# 0.06fF
C105 ffo_0/d xor_0/inv_1/op 0.52fF
C106 ffo_0/nand_0/b vdd 0.15fF
C107 ffo_0/nand_0/b ffo_0/nand_0/w_0_0# 0.06fF
C108 vdd ffo_0/inv_0/w_0_6# 0.06fF
C109 xor_0/inv_0/op k 0.27fF
C110 xor_0/inv_1/op vdd 0.15fF
C111 xor_0/w_n3_4# xor_0/inv_0/op 0.06fF
C112 vdd sbar 0.28fF
C113 ffo_0/nand_1/b gnd 0.26fF
C114 xor_0/a_10_10# Gnd 0.01fF
C115 xor_0/w_n3_4# Gnd 1.14fF
C116 xor_0/inv_1/op Gnd 0.49fF
C117 c Gnd 1.38fF
C118 xor_0/inv_1/w_0_6# Gnd 0.58fF
C119 xor_0/inv_0/op Gnd 0.50fF
C120 k Gnd 1.29fF
C121 xor_0/inv_0/w_0_6# Gnd 0.58fF
C122 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C123 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C124 gnd Gnd 3.20fF
C125 ffo_0/nand_7/a Gnd 0.30fF
C126 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C127 sbar Gnd 0.43fF
C128 vdd Gnd 1.79fF
C129 ffo_0/nand_6/a Gnd 0.30fF
C130 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C131 clk Gnd 1.06fF
C132 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C133 ffo_0/nand_3/b Gnd 0.43fF
C134 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C135 ffo_0/nand_3/a Gnd 0.30fF
C136 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C137 ffo_0/nand_0/b Gnd 0.63fF
C138 ffo_0/d Gnd 0.64fF
C139 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C140 ffo_0/inv_0/op Gnd 0.26fF
C141 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C142 ffo_0/nand_1/a Gnd 0.30fF
C143 ffo_0/nand_1/w_0_0# Gnd 0.82fF
