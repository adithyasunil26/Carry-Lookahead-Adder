magic
tech scmos
timestamp 1618500037
<< nwell >>
rect -6 2 46 38
<< ntransistor >>
rect 5 -32 7 -20
rect 12 -32 14 -20
rect 26 -32 28 -20
rect 33 -32 35 -20
<< ptransistor >>
rect 5 8 7 32
rect 12 8 14 32
rect 26 8 28 32
rect 33 8 35 32
<< ndiffusion >>
rect 0 -28 5 -20
rect 4 -32 5 -28
rect 7 -32 12 -20
rect 14 -24 18 -20
rect 22 -24 26 -20
rect 14 -32 26 -24
rect 28 -32 33 -20
rect 35 -28 40 -20
rect 35 -32 36 -28
<< pdiffusion >>
rect 4 28 5 32
rect 0 8 5 28
rect 7 8 12 32
rect 14 12 26 32
rect 14 8 18 12
rect 22 8 26 12
rect 28 8 33 32
rect 35 28 36 32
rect 35 8 40 28
<< ndcontact >>
rect 0 -32 4 -28
rect 18 -24 22 -20
rect 36 -32 40 -28
<< pdcontact >>
rect 0 28 4 32
rect 18 8 22 12
rect 36 28 40 32
<< polysilicon >>
rect 5 32 7 35
rect 12 32 14 35
rect 26 32 28 35
rect 33 32 35 35
rect 5 -20 7 8
rect 12 7 14 8
rect 26 7 28 8
rect 12 -20 14 -19
rect 26 -20 28 -19
rect 33 -20 35 8
rect 5 -35 7 -32
rect 12 -35 14 -32
rect 26 -35 28 -32
rect 33 -35 35 -32
<< polycontact >>
rect 1 -12 5 -8
rect 11 3 15 7
rect 25 3 29 7
rect 29 -5 33 -1
rect 11 -19 15 -15
rect 25 -19 29 -15
<< metal1 >>
rect -15 38 46 41
rect 0 32 3 38
rect 37 32 40 38
rect -51 10 -50 13
rect -15 10 -10 15
rect 19 -8 22 8
rect 19 -11 46 -8
rect -51 -21 -50 -18
rect -15 -22 -12 -18
rect 19 -20 22 -11
rect 0 -36 3 -32
rect 37 -36 40 -32
rect -6 -39 46 -36
<< m2contact >>
rect -50 9 -45 14
rect -50 -22 -45 -17
<< metal2 >>
rect -15 10 -10 15
rect -49 1 -46 9
rect 25 3 29 7
rect 25 1 28 3
rect -49 -2 -10 1
rect -13 -8 -10 -2
rect 12 -2 28 1
rect 12 -6 15 -2
rect -13 -11 5 -8
rect -48 -14 -17 -11
rect 1 -12 5 -11
rect 12 -9 22 -6
rect -48 -17 -45 -14
rect -20 -15 -17 -14
rect 12 -15 15 -9
rect -20 -16 -3 -15
rect 11 -16 15 -15
rect -20 -18 15 -16
rect -6 -19 15 -18
<< m123contact >>
rect -15 -27 -10 -22
<< metal3 >>
rect 11 3 15 7
rect 12 -5 15 3
rect -6 -6 15 -5
rect -6 -8 28 -6
rect -6 -23 -3 -8
rect 12 -9 28 -8
rect 25 -15 28 -9
rect 25 -19 29 -15
rect -10 -26 -3 -23
<< metal4 >>
rect -13 -2 -10 10
rect 29 -2 33 -1
rect -13 -5 33 -2
<< m345contact >>
rect -15 10 -10 15
use inv  inv_0
timestamp 1618367270
transform 1 0 -42 0 1 8
box -3 -13 27 33
use inv  inv_1
timestamp 1618367270
transform 1 0 -42 0 -1 -15
box -3 -13 27 33
<< labels >>
rlabel metal1 -51 -21 -51 -18 3 b
rlabel metal1 -51 10 -51 13 3 a
rlabel metal1 21 -38 21 -38 1 gnd!
rlabel metal1 46 -11 46 -8 7 op
rlabel metal1 20 40 20 40 5 vdd!
<< end >>
