* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 vdd a_39_n5# a_34_8# w_n3_2# pfet w=24 l=2
+  ad=0 pd=0 as=144 ps=60
M1005 a_34_n33# a_31_n20# op Gnd nfet w=12 l=2
+  ad=72 pd=36 as=168 ps=52
M1006 a_10_8# a_5_n13# vdd w_n3_2# pfet w=24 l=2
+  ad=144 pd=60 as=0 ps=0
M1007 a_10_n33# a_5_n13# gnd Gnd nfet w=12 l=2
+  ad=72 pd=36 as=0 ps=0
M1008 gnd a_39_n5# a_34_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 op a_14_2# a_10_8# w_n3_2# pfet w=24 l=2
+  ad=336 pd=76 as=0 ps=0
M1010 op a_14_n20# a_10_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_34_8# a_30_2# op w_n3_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd w_n3_2# 0.14fF
C1 inv_0/op gnd 0.10fF
C2 m3_n10_n50# b 0.03fF
C3 m2_n10_36# m3_n10_n50# 0.01fF
C4 op inv_1/op 0.19fF
C5 m2_n10_n50# m3_n10_n50# 0.01fF
C6 m2_39_n5# m3_n18_10# 0.02fF
C7 m3_n18_10# a_39_n5# 0.01fF
C8 m2_n10_36# vdd 0.04fF
C9 a_39_n5# a_30_2# 0.04fF
C10 m2_n10_n50# vdd 0.02fF
C11 a gnd 0.54fF
C12 w_n3_2# a_30_2# 0.08fF
C13 a_5_n13# a_14_2# 0.04fF
C14 inv_1/w_0_6# inv_1/op 0.03fF
C15 m3_n18_10# b 0.04fF
C16 b a_30_2# 0.03fF
C17 op gnd 0.04fF
C18 m3_n18_10# a_5_n13# 0.00fF
C19 m3_n10_n50# vdd 0.07fF
C20 inv_1/in inv_1/op 0.04fF
C21 b a 0.06fF
C22 op a_39_n5# 0.06fF
C23 op w_n3_2# 0.02fF
C24 m3_n10_n50# m3_n18_10# 0.07fF
C25 op b 0.21fF
C26 a a_5_n13# 0.04fF
C27 inv_0/w_0_6# vdd 0.06fF
C28 inv_1/in gnd 0.05fF
C29 vdd inv_0/op 0.15fF
C30 m1_39_n5# m2_39_n5# 0.01fF
C31 m1_39_n5# a_39_n5# 0.04fF
C32 m3_n10_n50# a 0.03fF
C33 m3_n18_10# inv_0/op 0.02fF
C34 inv_0/w_0_6# inv_0/op 0.03fF
C35 a vdd 0.02fF
C36 b inv_1/in 0.05fF
C37 a_31_n20# inv_1/op 0.03fF
C38 op vdd 0.03fF
C39 m3_n18_10# a 0.04fF
C40 inv_0/w_0_6# a 0.06fF
C41 a inv_0/op 0.04fF
C42 inv_1/op gnd 0.29fF
C43 vdd inv_1/w_0_6# 0.06fF
C44 op m3_n18_10# 0.01fF
C45 a_14_n20# b 0.03fF
C46 inv_1/op w_n3_2# 0.08fF
C47 vdd inv_1/in 0.02fF
C48 m1_39_n5# m3_n18_10# 0.00fF
C49 a_31_n20# a_39_n5# 0.04fF
C50 b inv_1/op 0.40fF
C51 a_14_n20# a_5_n13# 0.04fF
C52 inv_1/op a_5_n13# 0.00fF
C53 b gnd 0.16fF
C54 m2_39_n5# a_39_n5# 0.00fF
C55 m3_n10_n50# inv_1/op 0.04fF
C56 a_39_n5# w_n3_2# 0.06fF
C57 a inv_1/in 0.01fF
C58 inv_1/op a_14_2# 0.03fF
C59 op m1_39_n5# 0.07fF
C60 vdd inv_1/op 0.15fF
C61 m2_39_n5# b 0.01fF
C62 b w_n3_2# 0.08fF
C63 m3_n10_n50# gnd 0.01fF
C64 m3_n18_10# inv_1/op 0.25fF
C65 w_n3_2# a_5_n13# 0.06fF
C66 inv_1/w_0_6# inv_1/in 0.06fF
C67 b a_5_n13# 0.00fF
C68 m2_n18_10# m3_n18_10# 0.02fF
C69 m3_n18_10# gnd 0.01fF
C70 a inv_1/op 0.16fF
C71 m2_n18_10# inv_0/op 0.02fF
C72 w_n3_2# a_14_2# 0.08fF
C73 m3_n18_10# Gnd 0.07fF **FLOATING
C74 m3_n10_n50# Gnd 0.37fF **FLOATING
C75 m2_n10_n50# Gnd 0.09fF **FLOATING
C76 m2_39_n5# Gnd 0.08fF **FLOATING
C77 m2_n18_10# Gnd 0.09fF **FLOATING
C78 m2_n10_36# Gnd 0.07fF **FLOATING
C79 m1_39_n5# Gnd 0.02fF **FLOATING
C80 b Gnd 0.89fF **FLOATING
C81 a_31_n20# Gnd 0.09fF
C82 a_14_n20# Gnd 0.09fF
C83 op Gnd 0.11fF
C84 a_39_n5# Gnd 0.19fF
C85 a_30_2# Gnd 0.01fF
C86 a_14_2# Gnd 0.01fF
C87 a_5_n13# Gnd 0.19fF
C88 w_n3_2# Gnd 1.05fF
C89 gnd Gnd 0.54fF
C90 inv_1/op Gnd 0.30fF
C91 inv_1/in Gnd 0.14fF
C92 inv_1/w_0_6# Gnd 0.58fF
C93 inv_0/op Gnd 0.08fF
C94 vdd Gnd 0.29fF
C95 a Gnd 0.98fF
C96 inv_0/w_0_6# Gnd 0.58fF
