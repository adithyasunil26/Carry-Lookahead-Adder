* SPICE3 file created from ffi.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=540 ps=316
M1001 vdd nand_1/b nand_3/b nand_1/w_0_0# pfet w=12 l=2
+  ad=1080 pd=612 as=96 ps=40
M1002 nand_3/b nand_1/a vdd nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 nand_3/b nand_1/b nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd clk nand_1/a nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_1/a inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_1/a clk nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd clk nand_3/a nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 nand_3/a d vdd nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 nand_3/a clk nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd nand_3/b nand_1/b nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 nand_1/b nand_3/a vdd nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 nand_1/b nand_3/b nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd inv_1/op nand_6/a nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 nand_6/a nand_3/b vdd nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 nand_6/a inv_1/op nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 nand_5/a_13_n26# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd nand_1/b nand_7/a nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 nand_7/a inv_1/op vdd nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 nand_7/a nand_1/b nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 nand_6/a_13_n26# nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1025 vdd qbar q nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1026 q nand_6/a vdd nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 q qbar nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1028 nand_7/a_13_n26# nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1029 vdd q qbar nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1030 qbar nand_7/a vdd nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 qbar q nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1032 inv_0/op d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1033 inv_0/op d vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1034 inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1035 inv_1/op clk vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 nand_1/b nand_3/b 0.32fF
C1 nand_3/b nand_1/w_0_0# 0.04fF
C2 vdd nand_1/a 0.30fF
C3 inv_1/op nand_4/w_0_0# 0.06fF
C4 qbar q 0.32fF
C5 vdd nand_3/b 0.39fF
C6 inv_0/w_0_6# inv_0/op 0.03fF
C7 vdd q 0.28fF
C8 inv_1/op d 0.01fF
C9 inv_1/w_0_6# inv_1/op 0.04fF
C10 nand_3/w_0_0# nand_3/a 0.06fF
C11 nand_3/b nand_1/a 0.00fF
C12 gnd nand_7/a 0.03fF
C13 inv_0/op d 0.04fF
C14 nand_3/a nand_2/w_0_0# 0.04fF
C15 nand_7/a nand_1/b 0.13fF
C16 nand_6/a inv_1/op 0.13fF
C17 inv_1/op clk 0.07fF
C18 qbar nand_7/a 0.00fF
C19 inv_0/op clk 0.32fF
C20 nand_7/a vdd 0.30fF
C21 gnd inv_1/op 0.22fF
C22 gnd inv_0/op 0.10fF
C23 nand_2/w_0_0# d 0.06fF
C24 qbar nand_7/w_0_0# 0.04fF
C25 nand_1/b inv_1/op 0.45fF
C26 inv_0/op nand_0/w_0_0# 0.06fF
C27 nand_7/a q 0.31fF
C28 nand_7/w_0_0# vdd 0.10fF
C29 nand_3/a clk 0.13fF
C30 inv_0/w_0_6# d 0.06fF
C31 vdd inv_1/op 1.63fF
C32 gnd nand_3/a 0.03fF
C33 inv_0/op vdd 0.17fF
C34 nand_2/w_0_0# clk 0.06fF
C35 nand_1/b nand_5/w_0_0# 0.06fF
C36 nand_7/w_0_0# q 0.06fF
C37 nand_6/a nand_4/w_0_0# 0.04fF
C38 inv_1/op nand_3/b 0.33fF
C39 vdd nand_5/w_0_0# 0.10fF
C40 nand_3/w_0_0# nand_1/b 0.04fF
C41 nand_6/w_0_0# nand_6/a 0.06fF
C42 d clk 0.64fF
C43 inv_1/w_0_6# clk 0.06fF
C44 vdd nand_3/a 0.30fF
C45 nand_3/w_0_0# vdd 0.11fF
C46 gnd d 0.19fF
C47 vdd nand_2/w_0_0# 0.10fF
C48 nand_7/a nand_7/w_0_0# 0.06fF
C49 nand_3/b nand_3/a 0.31fF
C50 nand_3/w_0_0# nand_3/b 0.06fF
C51 vdd nand_4/w_0_0# 0.10fF
C52 inv_0/w_0_6# vdd 0.06fF
C53 qbar nand_6/w_0_0# 0.06fF
C54 gnd nand_6/a 0.03fF
C55 gnd clk 0.73fF
C56 nand_6/w_0_0# vdd 0.10fF
C57 vdd d 0.04fF
C58 vdd inv_1/w_0_6# 0.06fF
C59 nand_0/w_0_0# clk 0.06fF
C60 nand_3/b nand_4/w_0_0# 0.06fF
C61 nand_7/a nand_5/w_0_0# 0.04fF
C62 qbar nand_6/a 0.31fF
C63 nand_6/w_0_0# q 0.04fF
C64 nand_6/a vdd 0.30fF
C65 gnd nand_1/b 0.26fF
C66 vdd clk 0.02fF
C67 gnd qbar 0.52fF
C68 nand_1/a clk 0.13fF
C69 gnd vdd 0.03fF
C70 nand_1/b nand_1/w_0_0# 0.06fF
C71 inv_1/op nand_5/w_0_0# 0.06fF
C72 nand_6/a q 0.00fF
C73 gnd nand_1/a 0.03fF
C74 vdd nand_0/w_0_0# 0.10fF
C75 vdd nand_1/b 0.31fF
C76 vdd nand_1/w_0_0# 0.10fF
C77 gnd nand_3/b 0.35fF
C78 nand_1/a nand_0/w_0_0# 0.04fF
C79 qbar vdd 0.28fF
C80 gnd q 0.34fF
C81 nand_1/b nand_1/a 0.31fF
C82 nand_1/w_0_0# nand_1/a 0.06fF
C83 inv_1/w_0_6# Gnd 0.58fF
C84 inv_0/w_0_6# Gnd 0.58fF
C85 gnd Gnd 1.75fF
C86 nand_7/a Gnd 0.30fF
C87 nand_7/w_0_0# Gnd 0.82fF
C88 q Gnd 0.42fF
C89 vdd Gnd 1.12fF
C90 nand_6/a Gnd 0.30fF
C91 nand_6/w_0_0# Gnd 0.82fF
C92 inv_1/op Gnd 0.89fF
C93 nand_5/w_0_0# Gnd 0.82fF
C94 nand_3/b Gnd 0.43fF
C95 nand_4/w_0_0# Gnd 0.82fF
C96 nand_3/a Gnd 0.30fF
C97 nand_3/w_0_0# Gnd 0.82fF
C98 clk Gnd 0.89fF
C99 d Gnd 0.45fF
C100 nand_2/w_0_0# Gnd 0.82fF
C101 inv_0/op Gnd 0.26fF
C102 nand_0/w_0_0# Gnd 0.82fF
C103 nand_1/a Gnd 0.30fF
C104 nand_1/w_0_0# Gnd 0.82fF
