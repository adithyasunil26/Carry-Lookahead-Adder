* SPICE3 file created from ckt.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 gnd ffi_0/q inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in ffi_0/q nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd ffi_0/q inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in ffi_0/q nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1067 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1068 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a gnd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1071 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1072 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op gnd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1074 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1075 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1076 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1078 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1079 gnd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1080 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a gnd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1083 gnd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1084 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b gnd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1086 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1087 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1088 sumffo_0/ffo_0/nand_7/a clk gnd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1090 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1091 gnd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1092 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a gnd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1095 gnd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1096 z1o sumffo_0/ffo_0/nand_7/a gnd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1098 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1099 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1101 sumffo_0/ffo_0/nand_0/b clk gnd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1102 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_0/xor_0/inv_1/op ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_0/xor_0/inv_1/op ffi_0/q gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 gnd ffi_0/q sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 sumffo_0/ffo_0/d ffi_0/q sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1115 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1116 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a gnd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1119 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1120 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op gnd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1122 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1123 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1124 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1127 gnd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1128 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a gnd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1130 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1131 gnd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1132 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b gnd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1134 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1135 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1136 sumffo_2/ffo_0/nand_7/a clk gnd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1139 gnd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1140 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a gnd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1143 gnd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1144 z3o sumffo_2/ffo_0/nand_7/a gnd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1146 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1147 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 sumffo_2/ffo_0/nand_0/b clk gnd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1153 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1154 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1155 sumffo_2/ffo_0/d ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1156 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1157 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1158 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1163 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1164 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a gnd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1166 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1167 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1168 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op gnd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1170 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1171 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1172 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a gnd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1179 gnd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1180 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b gnd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1183 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1184 sumffo_1/ffo_0/nand_7/a clk gnd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1186 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1187 gnd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1188 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a gnd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1190 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1191 gnd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1192 z2o sumffo_1/ffo_0/nand_7/a gnd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1194 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1195 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 sumffo_1/ffo_0/nand_0/b clk gnd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1211 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1212 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a gnd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1214 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op gnd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1219 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1220 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1223 gnd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1224 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a gnd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1226 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1227 gnd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1228 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b gnd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1230 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1231 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1232 sumffo_3/ffo_0/nand_7/a clk gnd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1235 gnd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1236 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a gnd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1238 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1239 gnd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1240 z4o sumffo_3/ffo_0/nand_7/a gnd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1245 sumffo_3/ffo_0/nand_0/b clk gnd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1246 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1247 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1248 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1249 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1250 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1251 sumffo_3/ffo_0/d ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1252 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1253 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1254 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1259 gnd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1260 ffo_0/nand_3/b ffo_0/nand_1/a gnd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1262 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1263 gnd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1264 ffo_0/nand_1/a ffo_0/inv_0/op gnd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1266 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1267 gnd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1268 ffo_0/nand_3/a ffo_0/d gnd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1270 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1271 gnd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1272 ffo_0/nand_1/b ffo_0/nand_3/a gnd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1274 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1275 gnd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1276 ffo_0/nand_6/a ffo_0/nand_3/b gnd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1278 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1279 gnd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1280 ffo_0/nand_7/a clk gnd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1282 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1283 gnd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1284 ffo_0/qbar ffo_0/nand_6/a gnd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1286 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1287 gnd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1288 couto ffo_0/nand_7/a gnd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffo_0/inv_0/op ffo_0/d gnd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1293 ffo_0/nand_0/b clk gnd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1294 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1295 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1297 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1298 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1299 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1301 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1303 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1305 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1306 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1307 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1309 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1311 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1313 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1314 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1315 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1317 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1318 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1319 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1320 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1321 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1323 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1325 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1327 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1329 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1330 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1331 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipg_0/pggen_0/nand_0/a_13_n26# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 gnd ffipg_0/ffi_0/q cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 cla_0/g0 ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 cla_0/g0 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1337 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1338 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1339 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 gnd ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1341 ffipg_0/k ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1342 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1343 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1344 ffipg_0/pggen_0/xor_0/a_10_n43# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 nor_0/a ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1349 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 gnd ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1351 nor_0/a ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 ffipg_0/ffi_0/nand_1/a_13_n26# ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/a gnd ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipg_0/ffi_0/nand_0/a_13_n26# ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 gnd clk ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/inv_0/op gnd ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 ffipg_0/ffi_0/nand_1/a clk ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1361 gnd clk ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1362 ffipg_0/ffi_0/nand_3/a y1in gnd ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 ffipg_0/ffi_0/nand_3/a clk ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipg_0/ffi_0/nand_3/a_13_n26# ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 gnd ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/a gnd ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipg_0/ffi_0/nand_4/a_13_n26# ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1369 gnd ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1370 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_3/b gnd ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1371 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 ffipg_0/ffi_0/nand_5/a_13_n26# ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1373 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1374 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/inv_1/op gnd ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1376 ffipg_0/ffi_0/nand_6/a_13_n26# ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1377 gnd ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1378 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/a gnd ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1380 ffipg_0/ffi_0/nand_7/a_13_n26# ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1381 gnd ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1382 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a gnd ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1384 ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1385 ffipg_0/ffi_0/inv_0/op y1in gnd ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1386 ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1387 ffipg_0/ffi_0/inv_1/op clk gnd ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipg_0/ffi_1/nand_1/a_13_n26# ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a gnd ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipg_0/ffi_1/nand_0/a_13_n26# ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 gnd clk ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/inv_0/op gnd ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipg_0/ffi_1/nand_1/a clk ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 gnd clk ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipg_0/ffi_1/nand_3/a x1in gnd ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipg_0/ffi_1/nand_3/a clk ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipg_0/ffi_1/nand_3/a_13_n26# ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 gnd ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/a gnd ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipg_0/ffi_1/nand_4/a_13_n26# ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 gnd ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_3/b gnd ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipg_0/ffi_1/nand_5/a_13_n26# ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/inv_1/op gnd ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipg_0/ffi_1/nand_6/a_13_n26# ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 gnd ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/a gnd ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipg_0/ffi_1/nand_7/a_13_n26# ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1417 gnd ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1418 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a gnd ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1421 ffipg_0/ffi_1/inv_0/op x1in gnd ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1422 ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1423 ffipg_0/ffi_1/inv_1/op clk gnd ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1425 ffo_0/d inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1426 ffipg_1/pggen_0/nand_0/a_13_n26# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1427 gnd ffipg_1/ffi_0/q cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 cla_0/l ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 cla_0/l ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1431 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1433 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1434 gnd ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1435 ffipg_1/k ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1436 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1437 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1438 ffipg_1/pggen_0/xor_0/a_10_n43# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 cla_1/p0 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1443 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 gnd ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1445 cla_1/p0 ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 ffipg_1/ffi_0/nand_1/a_13_n26# ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1447 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1448 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a gnd ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1450 ffipg_1/ffi_0/nand_0/a_13_n26# ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1451 gnd clk ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1452 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/inv_0/op gnd ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 ffipg_1/ffi_0/nand_1/a clk ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1455 gnd clk ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1456 ffipg_1/ffi_0/nand_3/a y2in gnd ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 ffipg_1/ffi_0/nand_3/a clk ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1458 ffipg_1/ffi_0/nand_3/a_13_n26# ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1459 gnd ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1460 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/a gnd ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 ffipg_1/ffi_0/nand_4/a_13_n26# ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1463 gnd ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1464 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_3/b gnd ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1466 ffipg_1/ffi_0/nand_5/a_13_n26# ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1467 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1468 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/inv_1/op gnd ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1470 ffipg_1/ffi_0/nand_6/a_13_n26# ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 gnd ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a gnd ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 ffipg_1/ffi_0/nand_7/a_13_n26# ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 gnd ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a gnd ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 ffipg_1/ffi_0/inv_0/op y2in gnd ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1480 ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1481 ffipg_1/ffi_0/inv_1/op clk gnd ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 ffipg_1/ffi_1/nand_1/a_13_n26# ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a gnd ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 ffipg_1/ffi_1/nand_0/a_13_n26# ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 gnd clk ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/inv_0/op gnd ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 ffipg_1/ffi_1/nand_1/a clk ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 gnd clk ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 ffipg_1/ffi_1/nand_3/a x2in gnd ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 ffipg_1/ffi_1/nand_3/a clk ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 ffipg_1/ffi_1/nand_3/a_13_n26# ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 gnd ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/a gnd ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 ffipg_1/ffi_1/nand_4/a_13_n26# ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 gnd ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_3/b gnd ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 ffipg_1/ffi_1/nand_5/a_13_n26# ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1503 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1504 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/inv_1/op gnd ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1505 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 ffipg_1/ffi_1/nand_6/a_13_n26# ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1507 gnd ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1508 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a gnd ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 ffipg_1/ffi_1/nand_7/a_13_n26# ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1511 gnd ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1512 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a gnd ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1513 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1514 ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1515 ffipg_1/ffi_1/inv_0/op x2in gnd ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1516 ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1517 ffipg_1/ffi_1/inv_1/op clk gnd ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1518 ffipg_2/pggen_0/nand_0/a_13_n26# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 gnd ffipg_2/ffi_0/q cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1520 cla_0/l ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 cla_0/l ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1523 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1524 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1525 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 gnd ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1527 ffipg_2/k ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1528 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1529 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1530 ffipg_2/pggen_0/xor_0/a_10_n43# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1534 cla_2/p0 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1535 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 gnd ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1537 cla_2/p0 ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 ffipg_2/ffi_0/nand_1/a_13_n26# ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a gnd ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 ffipg_2/ffi_0/nand_0/a_13_n26# ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 gnd clk ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/inv_0/op gnd ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 ffipg_2/ffi_0/nand_1/a clk ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 gnd clk ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 ffipg_2/ffi_0/nand_3/a y3in gnd ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 ffipg_2/ffi_0/nand_3/a clk ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 ffipg_2/ffi_0/nand_3/a_13_n26# ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1551 gnd ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1552 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/a gnd ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 ffipg_2/ffi_0/nand_4/a_13_n26# ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1555 gnd ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1556 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_3/b gnd ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 ffipg_2/ffi_0/nand_5/a_13_n26# ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1559 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1560 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/inv_1/op gnd ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1561 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1562 ffipg_2/ffi_0/nand_6/a_13_n26# ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1563 gnd ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1564 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/a gnd ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1566 ffipg_2/ffi_0/nand_7/a_13_n26# ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 gnd ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a gnd ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1571 ffipg_2/ffi_0/inv_0/op y3in gnd ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1572 ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1573 ffipg_2/ffi_0/inv_1/op clk gnd ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 ffipg_2/ffi_1/nand_1/a_13_n26# ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a gnd ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 ffipg_2/ffi_1/nand_0/a_13_n26# ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 gnd clk ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/inv_0/op gnd ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 ffipg_2/ffi_1/nand_1/a clk ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 gnd clk ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 ffipg_2/ffi_1/nand_3/a x3in gnd ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 ffipg_2/ffi_1/nand_3/a clk ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 ffipg_2/ffi_1/nand_3/a_13_n26# ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 gnd ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/a gnd ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 ffipg_2/ffi_1/nand_4/a_13_n26# ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 gnd ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_3/b gnd ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 ffipg_2/ffi_1/nand_5/a_13_n26# ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/inv_1/op gnd ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 ffipg_2/ffi_1/nand_6/a_13_n26# ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1599 gnd ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1600 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/a gnd ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1601 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 ffipg_2/ffi_1/nand_7/a_13_n26# ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1603 gnd ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1604 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a gnd ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1605 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1607 ffipg_2/ffi_1/inv_0/op x3in gnd ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1608 ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1609 ffipg_2/ffi_1/inv_1/op clk gnd ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1610 ffi_0/nand_1/a_13_n26# ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1611 gnd ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1612 ffi_0/nand_3/b ffi_0/nand_1/a gnd ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1614 ffi_0/nand_0/a_13_n26# ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 gnd clk ffi_0/nand_1/a ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 ffi_0/nand_1/a ffi_0/inv_0/op gnd ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 ffi_0/nand_1/a clk ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 gnd clk ffi_0/nand_3/a ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 ffi_0/nand_3/a cinin gnd ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 ffi_0/nand_3/a clk ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 ffi_0/nand_3/a_13_n26# ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 gnd ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 ffi_0/nand_1/b ffi_0/nand_3/a gnd ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 ffi_0/nand_4/a_13_n26# ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 gnd ffi_0/inv_1/op ffi_0/nand_6/a ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 ffi_0/nand_6/a ffi_0/nand_3/b gnd ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 ffi_0/nand_6/a ffi_0/inv_1/op ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 ffi_0/nand_5/a_13_n26# ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 gnd ffi_0/nand_1/b ffi_0/nand_7/a ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 ffi_0/nand_7/a ffi_0/inv_1/op gnd ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 ffi_0/nand_7/a ffi_0/nand_1/b ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 ffi_0/nand_6/a_13_n26# ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 gnd ffi_0/q nor_0/b ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 nor_0/b ffi_0/nand_6/a gnd ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 nor_0/b ffi_0/q ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 ffi_0/nand_7/a_13_n26# ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 gnd nor_0/b ffi_0/q ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 ffi_0/q ffi_0/nand_7/a gnd ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 ffi_0/q nor_0/b ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1643 ffi_0/inv_0/op cinin gnd ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1644 ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1645 ffi_0/inv_1/op clk gnd ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 ffipg_3/pggen_0/nand_0/a_13_n26# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1647 gnd ffipg_3/ffi_0/q cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1648 cla_2/g1 ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1649 cla_2/g1 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 gnd ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 ffipg_3/k ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 ffipg_3/pggen_0/xor_0/a_10_n43# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 cla_2/p1 ffipg_3/ffi_1/q ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1663 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 gnd ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1665 cla_2/p1 ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1666 ffipg_3/ffi_0/nand_1/a_13_n26# ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/a gnd ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffipg_3/ffi_0/nand_0/a_13_n26# ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 gnd clk ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/inv_0/op gnd ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffipg_3/ffi_0/nand_1/a clk ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 gnd clk ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffipg_3/ffi_0/nand_3/a y4in gnd ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffipg_3/ffi_0/nand_3/a clk ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffipg_3/ffi_0/nand_3/a_13_n26# ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 gnd ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/a gnd ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffipg_3/ffi_0/nand_4/a_13_n26# ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 gnd ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_3/b gnd ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffipg_3/ffi_0/nand_5/a_13_n26# ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/inv_1/op gnd ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffipg_3/ffi_0/nand_6/a_13_n26# ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 gnd ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/a gnd ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffipg_3/ffi_0/nand_7/a_13_n26# ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1695 gnd ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1696 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a gnd ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1697 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 ffipg_3/ffi_0/inv_0/op y4in gnd ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 ffipg_3/ffi_0/inv_1/op clk gnd ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 ffipg_3/ffi_1/nand_1/a_13_n26# ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1703 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1704 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/a gnd ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1705 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1706 ffipg_3/ffi_1/nand_0/a_13_n26# ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1707 gnd clk ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1708 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/inv_0/op gnd ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1709 ffipg_3/ffi_1/nand_1/a clk ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1711 gnd clk ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1712 ffipg_3/ffi_1/nand_3/a x4in gnd ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1713 ffipg_3/ffi_1/nand_3/a clk ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1714 ffipg_3/ffi_1/nand_3/a_13_n26# ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1715 gnd ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1716 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/a gnd ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1717 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1718 ffipg_3/ffi_1/nand_4/a_13_n26# ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1719 gnd ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1720 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_3/b gnd ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1721 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 ffipg_3/ffi_1/nand_5/a_13_n26# ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1723 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1724 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/inv_1/op gnd ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1725 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1726 ffipg_3/ffi_1/nand_6/a_13_n26# ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1727 gnd ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1728 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/a gnd ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1730 ffipg_3/ffi_1/nand_7/a_13_n26# ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1731 gnd ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1732 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a gnd ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 ffipg_3/ffi_1/inv_0/op x4in gnd ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffipg_3/ffi_1/inv_1/op clk gnd ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 cla_2/inv_0/in cla_2/p1 0.02fF
C1 gnd ffipg_2/ffi_1/nand_0/a_13_n26# 0.01fF
C2 sumffo_1/ffo_0/d clk 0.04fF
C3 ffi_0/nand_6/a ffi_0/q 0.31fF
C4 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/inv_1/op 0.33fF
C5 sumffo_3/xor_0/w_n3_4# ffipg_3/k 0.06fF
C6 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C7 ffo_0/nand_6/a clk 0.13fF
C8 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/sbar 0.04fF
C9 ffipg_0/ffi_0/nand_1/a gnd 0.44fF
C10 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C11 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# 0.04fF
C12 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C13 inv_8/in ffi_0/q 0.13fF
C14 nor_4/a inv_9/in 0.02fF
C15 gnd ffipg_3/ffi_1/inv_0/op 0.27fF
C16 gnd ffipg_3/ffi_0/nand_1/w_0_0# 0.10fF
C17 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/inv_1/op 0.33fF
C18 ffipg_0/ffi_0/nand_0/w_0_0# ffipg_0/ffi_0/inv_0/op 0.06fF
C19 sumffo_0/sbar sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C20 ffipg_0/ffi_0/nand_0/w_0_0# clk 0.06fF
C21 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C22 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C23 gnd nor_2/w_0_0# 0.15fF
C24 sumffo_1/ffo_0/nand_6/a sumffo_1/sbar 0.00fF
C25 sumffo_0/ffo_0/nand_3/b gnd 0.74fF
C26 ffipg_2/ffi_0/inv_0/w_0_6# y3in 0.06fF
C27 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C28 inv_8/w_0_6# ffi_0/q 0.06fF
C29 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C30 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C31 sumffo_0/ffo_0/nand_0/a_13_n26# gnd 0.01fF
C32 gnd ffipg_2/ffi_1/nand_5/w_0_0# 0.10fF
C33 gnd ffipg_3/ffi_0/nand_0/w_0_0# 0.10fF
C34 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C35 ffipg_2/ffi_0/nand_6/a gnd 0.37fF
C36 gnd ffipg_3/ffi_1/nand_0/w_0_0# 0.10fF
C37 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/b 0.31fF
C38 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar 0.32fF
C39 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/inv_1/w_0_6# 0.04fF
C40 ffipg_0/k ffi_0/q 0.19fF
C41 inv_6/in nor_3/w_0_0# 0.11fF
C42 gnd ffipg_3/ffi_1/nand_3/a 0.33fF
C43 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C44 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b 0.13fF
C45 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_3/b 0.00fF
C46 ffipg_1/ffi_0/inv_0/op y2in 0.04fF
C47 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C48 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C49 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C50 inv_4/in cla_1/n 0.02fF
C51 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# 0.04fF
C52 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C53 cla_1/inv_0/op cla_0/l 0.35fF
C54 ffipg_2/ffi_0/nand_1/w_0_0# gnd 0.10fF
C55 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_3/b 0.04fF
C56 inv_0/op cla_0/g0 0.33fF
C57 sumffo_3/xor_0/a_10_10# ffi_0/q 0.04fF
C58 x4in ffipg_3/ffi_1/inv_1/op 0.01fF
C59 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C60 ffipg_1/ffi_0/nand_1/a clk 0.13fF
C61 nand_2/b cla_0/n 0.06fF
C62 ffipg_1/ffi_1/nand_3/a clk 0.13fF
C63 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a 0.31fF
C64 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_7/a 0.04fF
C65 cla_2/l inv_7/w_0_6# 0.06fF
C66 clk ffipg_3/ffi_0/inv_1/op 0.07fF
C67 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C68 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C69 gnd ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C70 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_1/b 0.45fF
C71 inv_5/in nor_3/b 0.04fF
C72 ffo_0/nand_3/b ffo_0/nand_3/w_0_0# 0.06fF
C73 gnd inv_3/in 0.47fF
C74 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C75 gnd z1o 0.80fF
C76 gnd ffipg_1/ffi_1/nand_3/w_0_0# 0.11fF
C77 gnd ffipg_0/ffi_1/qbar 0.67fF
C78 cla_2/l cla_2/p1 0.02fF
C79 cla_2/l cla_0/n 0.32fF
C80 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/inv_1/w_0_6# 0.04fF
C81 ffo_0/nand_6/a couto 0.31fF
C82 ffipg_0/ffi_1/nand_2/w_0_0# x1in 0.06fF
C83 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_1/q 0.06fF
C84 ffipg_2/pggen_0/nand_0/w_0_0# ffipg_2/ffi_0/q 0.06fF
C85 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C86 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a 0.00fF
C87 gnd ffipg_2/ffi_0/nand_7/w_0_0# 0.10fF
C88 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C89 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/ffi_0/q 0.23fF
C90 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q 0.27fF
C91 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C92 sumffo_1/ffo_0/nand_6/w_0_0# gnd 0.10fF
C93 cla_0/inv_0/in cla_0/l 0.07fF
C94 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C95 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/inv_1/op 0.45fF
C96 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_0/b 0.06fF
C97 gnd ffipg_3/ffi_0/nand_4/w_0_0# 0.10fF
C98 gnd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C99 ffipg_1/ffi_1/inv_1/op x2in 0.01fF
C100 ffo_0/nand_7/w_0_0# couto 0.04fF
C101 sumffo_0/ffo_0/nand_6/a clk 0.13fF
C102 gnd cla_2/nand_0/a_13_n26# 0.01fF
C103 y2in ffipg_1/ffi_0/inv_1/op 0.01fF
C104 nor_1/b inv_2/w_0_6# 0.03fF
C105 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C106 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C107 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/inv_0/w_0_6# 0.03fF
C108 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C109 ffipg_1/ffi_1/inv_0/op clk 0.32fF
C110 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/q 0.31fF
C111 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/qbar 0.04fF
C112 gnd ffipg_0/ffi_0/nand_5/w_0_0# 0.10fF
C113 sumffo_1/ffo_0/nand_6/a gnd 0.33fF
C114 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# 0.04fF
C115 sumffo_2/ffo_0/nand_3/b clk 0.33fF
C116 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C117 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_1/b 0.31fF
C118 gnd ffipg_0/ffi_1/nand_3/b 0.74fF
C119 y4in ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C120 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/nand_6/a 0.04fF
C121 gnd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C122 sumffo_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C123 cla_1/p0 nor_0/a 0.24fF
C124 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a 0.31fF
C125 gnd ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C126 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C127 gnd sumffo_1/ffo_0/nand_4/w_0_0# 0.10fF
C128 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/inv_1/op 0.33fF
C129 ffipg_0/pggen_0/nand_0/w_0_0# cla_0/g0 0.04fF
C130 ffipg_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C131 clk ffipg_3/ffi_0/nand_1/a 0.13fF
C132 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a 0.00fF
C133 gnd ffipg_0/ffi_1/nand_0/a_13_n26# 0.01fF
C134 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C135 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q 0.22fF
C136 gnd ffipg_1/ffi_0/nand_7/a 0.37fF
C137 sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d 0.06fF
C138 gnd cla_2/inv_0/in 0.34fF
C139 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C140 ffipg_3/ffi_1/nand_0/w_0_0# ffipg_3/ffi_1/inv_0/op 0.06fF
C141 inv_4/in nor_2/b 0.16fF
C142 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/b 0.31fF
C143 sumffo_3/xor_0/w_n3_4# gnd 0.12fF
C144 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C145 cla_0/l ffipg_1/ffi_0/q 0.13fF
C146 gnd ffipg_3/ffi_1/nand_7/w_0_0# 0.10fF
C147 ffi_0/nand_7/w_0_0# ffi_0/q 0.04fF
C148 sumffo_2/ffo_0/nand_0/b clk 0.04fF
C149 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C150 gnd ffi_0/q 2.14fF
C151 sumffo_3/ffo_0/nand_1/w_0_0# gnd 0.10fF
C152 ffo_0/d nor_4/w_0_0# 0.03fF
C153 gnd sumffo_0/ffo_0/nand_1/b 0.57fF
C154 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/qbar 0.31fF
C155 gnd ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C156 sumffo_3/xor_0/a_38_n43# ffi_0/q 0.01fF
C157 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C158 sumffo_3/ffo_0/nand_5/w_0_0# clk 0.06fF
C159 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C160 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C161 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C162 sumffo_0/ffo_0/d gnd 0.41fF
C163 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/nand_7/a 0.04fF
C164 inv_1/in nor_1/w_0_0# 0.11fF
C165 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/op 0.04fF
C166 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C167 inv_0/in gnd 0.30fF
C168 ffipg_0/k nor_0/a 0.05fF
C169 gnd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C170 ffipg_1/ffi_0/nand_2/w_0_0# clk 0.06fF
C171 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C172 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C173 ffipg_2/ffi_1/inv_0/op clk 0.32fF
C174 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_1/b 0.04fF
C175 inv_2/in nor_1/b 0.04fF
C176 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C177 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C178 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_1/a 0.06fF
C179 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.35fF
C180 sumffo_1/ffo_0/nand_0/b clk 0.04fF
C181 gnd sumffo_0/ffo_0/nand_0/w_0_0# 0.10fF
C182 cla_2/nor_1/w_0_0# gnd 0.31fF
C183 ffipg_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C184 ffipg_1/k cla_0/g0 0.06fF
C185 nand_2/b gnd 1.90fF
C186 sumffo_1/xor_0/a_10_10# ffi_0/q 0.04fF
C187 gnd ffipg_2/ffi_1/inv_1/op 1.85fF
C188 gnd ffipg_1/ffi_0/nand_6/a 0.37fF
C189 gnd ffipg_1/ffi_1/nand_6/a 0.37fF
C190 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/inv_1/op 0.06fF
C191 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C192 inv_3/w_0_6# nor_2/b 0.03fF
C193 gnd ffipg_1/ffi_1/nand_1/b 0.57fF
C194 ffo_0/nand_3/b ffo_0/nand_4/w_0_0# 0.06fF
C195 gnd sumffo_0/ffo_0/nand_2/w_0_0# 0.10fF
C196 gnd cla_2/l 0.58fF
C197 ffipg_2/ffi_0/nand_3/w_0_0# gnd 0.11fF
C198 ffipg_0/pggen_0/nand_0/w_0_0# ffipg_0/ffi_0/q 0.06fF
C199 ffi_0/nand_3/a ffi_0/nand_3/w_0_0# 0.06fF
C200 nor_0/w_0_0# ffi_0/q 0.16fF
C201 ffipg_1/pggen_0/nor_0/w_0_0# cla_1/p0 0.05fF
C202 y2in ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C203 y1in ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C204 inv_1/in cla_0/n 0.02fF
C205 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C206 sumffo_1/ffo_0/nand_3/w_0_0# gnd 0.11fF
C207 clk ffipg_3/ffi_0/nand_3/a 0.13fF
C208 gnd cla_0/nor_0/w_0_0# 0.31fF
C209 ffo_0/nand_5/w_0_0# ffo_0/nand_7/a 0.04fF
C210 ffo_0/d gnd 0.45fF
C211 sumffo_1/xor_0/inv_1/op gnd 0.35fF
C212 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C213 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/nand_7/a 0.06fF
C214 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q 0.27fF
C215 nand_2/b ffipg_2/k 0.06fF
C216 gnd ffipg_1/ffi_1/nand_1/w_0_0# 0.10fF
C217 ffi_0/nand_4/w_0_0# ffi_0/nand_6/a 0.04fF
C218 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a 0.13fF
C219 gnd ffipg_2/ffi_1/q 2.24fF
C220 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# 0.04fF
C221 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C222 gnd cla_0/nand_0/w_0_0# 0.10fF
C223 sumffo_2/xor_0/a_10_10# gnd 0.93fF
C224 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_3/b 0.04fF
C225 gnd cla_2/n 0.60fF
C226 ffipg_2/ffi_1/nand_4/w_0_0# ffipg_2/ffi_1/inv_1/op 0.06fF
C227 cla_0/l ffipg_2/ffi_0/q 0.13fF
C228 ffipg_1/ffi_1/inv_0/op ffipg_1/ffi_1/nand_0/w_0_0# 0.06fF
C229 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C230 inv_0/in nor_0/w_0_0# 0.11fF
C231 ffo_0/inv_1/w_0_6# ffo_0/nand_0/b 0.03fF
C232 gnd ffipg_3/ffi_0/nand_7/w_0_0# 0.10fF
C233 gnd sumffo_3/ffo_0/nand_0/b 0.53fF
C234 sumffo_2/ffo_0/nand_6/a gnd 0.33fF
C235 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b 0.32fF
C236 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a 0.31fF
C237 gnd ffipg_3/ffi_1/qbar 0.67fF
C238 ffi_0/nand_7/w_0_0# ffi_0/nand_7/a 0.06fF
C239 gnd ffi_0/nand_7/a 0.33fF
C240 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C241 gnd ffipg_1/ffi_0/nand_0/w_0_0# 0.10fF
C242 gnd ffipg_0/ffi_0/inv_1/op 1.85fF
C243 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# 0.04fF
C244 clk ffipg_3/ffi_0/inv_0/op 0.32fF
C245 nor_1/b nor_1/w_0_0# 0.06fF
C246 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C247 gnd ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C248 inv_4/op inv_4/in 0.04fF
C249 sumffo_3/ffo_0/nand_3/b clk 0.33fF
C250 gnd sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C251 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a 0.00fF
C252 sumffo_1/ffo_0/nand_2/w_0_0# gnd 0.10fF
C253 gnd ffipg_3/ffi_0/nand_3/b 0.74fF
C254 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a 0.00fF
C255 gnd sumffo_3/ffo_0/nand_3/w_0_0# 0.11fF
C256 nand_2/b nor_0/w_0_0# 0.04fF
C257 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C258 ffipg_2/k ffipg_2/ffi_1/q 0.46fF
C259 ffo_0/nand_0/w_0_0# ffo_0/nand_0/b 0.06fF
C260 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar 0.32fF
C261 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/qbar 0.00fF
C262 ffi_0/nand_3/b ffi_0/nand_4/w_0_0# 0.06fF
C263 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C264 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C265 gnd nor_0/a 0.54fF
C266 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C267 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C268 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/ffi_1/q 0.06fF
C269 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/w_0_0# 0.06fF
C270 ffipg_2/ffi_0/inv_0/op clk 0.32fF
C271 gnd ffipg_2/ffi_0/qbar 0.67fF
C272 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/ffo_0/nand_6/a 0.06fF
C273 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C274 gnd sumffo_2/xor_0/inv_1/op 0.35fF
C275 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_1/w_0_6# 0.03fF
C276 ffipg_2/ffi_0/nand_2/w_0_0# clk 0.06fF
C277 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b 0.32fF
C278 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C279 inv_3/w_0_6# cla_0/n 0.16fF
C280 gnd ffipg_2/ffi_1/nand_6/w_0_0# 0.10fF
C281 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_1/b 0.06fF
C282 gnd ffipg_0/ffi_1/nand_1/a 0.45fF
C283 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# 0.04fF
C284 cinin clk 0.68fF
C285 gnd ffipg_3/ffi_1/nand_5/w_0_0# 0.10fF
C286 ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C287 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C288 ffipg_1/ffi_0/nand_3/w_0_0# ffipg_1/ffi_0/nand_3/b 0.06fF
C289 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/inv_1/op 0.06fF
C290 nor_1/b cla_0/n 0.36fF
C291 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b 0.32fF
C292 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C293 gnd ffo_0/inv_0/w_0_6# 0.07fF
C294 cla_1/l cla_0/l 0.08fF
C295 ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C296 gnd ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C297 gnd ffipg_3/ffi_1/nand_1/a 0.44fF
C298 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# 0.04fF
C299 ffipg_2/ffi_0/inv_0/op y3in 0.04fF
C300 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/qbar 0.00fF
C301 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.32fF
C302 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C303 y3in ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C304 gnd ffipg_0/ffi_0/nand_2/w_0_0# 0.10fF
C305 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/sbar 0.06fF
C306 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C307 ffipg_2/ffi_0/nand_3/b gnd 0.74fF
C308 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b 0.32fF
C309 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/ffi_0/q 0.12fF
C310 ffipg_0/pggen_0/nand_0/w_0_0# ffipg_0/ffi_1/q 0.06fF
C311 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C312 sumffo_2/ffo_0/nand_4/w_0_0# clk 0.06fF
C313 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C314 gnd ffo_0/qbar 0.62fF
C315 gnd ffo_0/nand_3/a 0.49fF
C316 gnd sumffo_0/xor_0/inv_1/op 0.35fF
C317 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_7/a 0.04fF
C318 nand_2/b inv_3/in 0.13fF
C319 sumffo_0/xor_0/inv_1/w_0_6# ffi_0/q 0.23fF
C320 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k 0.06fF
C321 gnd ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C322 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/a 0.06fF
C323 sumffo_2/ffo_0/nand_5/w_0_0# clk 0.06fF
C324 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_1/inv_1/op 0.75fF
C325 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b 0.32fF
C326 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C327 gnd ffipg_0/ffi_0/inv_0/op 0.27fF
C328 inv_1/in gnd 0.35fF
C329 sumffo_1/ffo_0/nand_3/b clk 0.33fF
C330 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_0/op 0.32fF
C331 gnd clk 24.51fF
C332 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C333 nor_0/w_0_0# nor_0/a 0.06fF
C334 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/q 0.06fF
C335 gnd inv_4/in 0.33fF
C336 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/ffi_0/q 0.06fF
C337 gnd ffipg_0/ffi_1/inv_1/op 1.85fF
C338 ffo_0/nand_2/w_0_0# gnd 0.10fF
C339 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# 0.04fF
C340 sumffo_3/xor_0/w_n3_4# ffi_0/q 0.01fF
C341 ffipg_2/ffi_1/nand_2/w_0_0# x3in 0.06fF
C342 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C343 ffipg_1/k ffipg_1/ffi_0/q 0.07fF
C344 cla_2/g1 cla_2/p1 0.00fF
C345 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_3/b 0.04fF
C346 gnd ffo_0/nand_1/b 0.57fF
C347 cla_1/inv_0/in cla_0/l 0.23fF
C348 gnd ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C349 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# 0.04fF
C350 gnd y1in 0.22fF
C351 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a 0.13fF
C352 ffipg_2/ffi_1/nand_3/a clk 0.13fF
C353 cla_2/p0 cla_1/p0 0.24fF
C354 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C355 ffi_0/nand_5/w_0_0# ffi_0/inv_1/op 0.06fF
C356 gnd ffi_0/nand_4/w_0_0# 0.10fF
C357 ffipg_1/pggen_0/nor_0/w_0_0# gnd 0.11fF
C358 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C359 gnd y3in 0.22fF
C360 gnd ffipg_0/ffi_1/nand_6/w_0_0# 0.10fF
C361 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_7/w_0_0# 0.06fF
C362 sumffo_2/xor_0/a_38_n43# ffi_0/q 0.01fF
C363 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# 0.04fF
C364 sumffo_3/ffo_0/nand_1/b clk 0.45fF
C365 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d 0.04fF
C366 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C367 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C368 cla_0/g0 cla_1/p0 0.38fF
C369 sumffo_1/ffo_0/nand_5/w_0_0# gnd 0.10fF
C370 sumffo_0/ffo_0/nand_4/w_0_0# gnd 0.10fF
C371 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a 0.00fF
C372 cla_2/p0 ffipg_3/k 0.06fF
C373 inv_0/in ffi_0/q 0.07fF
C374 ffi_0/nand_2/w_0_0# cinin 0.06fF
C375 gnd ffipg_0/ffi_1/nand_6/a 0.37fF
C376 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C377 cla_2/p0 cla_2/p1 0.24fF
C378 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/qbar 0.00fF
C379 gnd ffipg_1/ffi_1/nand_2/w_0_0# 0.10fF
C380 ffipg_3/ffi_0/nand_2/w_0_0# y4in 0.06fF
C381 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C382 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.32fF
C383 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C384 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C385 sumffo_1/ffo_0/nand_7/w_0_0# gnd 0.10fF
C386 sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# 0.04fF
C387 gnd cla_0/inv_0/op 0.27fF
C388 nand_2/b ffi_0/q 0.04fF
C389 ffi_0/inv_0/op ffi_0/nand_0/w_0_0# 0.06fF
C390 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C391 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# 0.04fF
C392 gnd couto 0.80fF
C393 gnd inv_3/w_0_6# 0.17fF
C394 sumffo_2/ffo_0/inv_1/w_0_6# sumffo_2/ffo_0/nand_0/b 0.03fF
C395 nor_4/w_0_0# inv_9/in 0.11fF
C396 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b 0.13fF
C397 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C398 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C399 gnd ffipg_3/ffi_1/nand_4/w_0_0# 0.10fF
C400 ffipg_0/ffi_0/nand_1/a clk 0.13fF
C401 gnd nor_1/b 0.35fF
C402 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C403 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.35fF
C404 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C405 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C406 gnd ffi_0/nand_2/w_0_0# 0.10fF
C407 sumffo_1/xor_0/inv_1/op ffi_0/q 0.04fF
C408 clk ffipg_3/ffi_1/inv_0/op 0.32fF
C409 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C410 cla_2/inv_0/op cla_2/g1 0.35fF
C411 gnd ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C412 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C413 gnd ffipg_1/ffi_0/nand_6/w_0_0# 0.10fF
C414 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C415 sumffo_0/ffo_0/nand_3/b clk 0.33fF
C416 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C417 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_0/b 0.40fF
C418 gnd ffipg_3/ffi_1/nand_2/w_0_0# 0.10fF
C419 inv_4/in nor_2/w_0_0# 0.11fF
C420 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/qbar 0.06fF
C421 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C422 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C423 gnd ffipg_2/ffi_1/nand_3/w_0_0# 0.11fF
C424 clk ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C425 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C426 sumffo_2/xor_0/a_10_10# ffi_0/q 0.04fF
C427 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C428 clk ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C429 ffipg_3/ffi_0/inv_0/op ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C430 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C431 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a 0.13fF
C432 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b 0.32fF
C433 sumffo_1/ffo_0/nand_1/b gnd 0.57fF
C434 gnd sumffo_0/ffo_0/nand_3/a 0.33fF
C435 gnd ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C436 sumffo_2/ffo_0/nand_1/w_0_0# gnd 0.10fF
C437 clk ffipg_3/ffi_1/nand_3/a 0.13fF
C438 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C439 gnd ffipg_3/ffi_1/nand_7/a 0.37fF
C440 ffi_0/nand_7/a ffi_0/q 0.00fF
C441 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C442 ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.32fF
C443 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/a 0.06fF
C444 gnd nor_3/b 0.33fF
C445 sumffo_1/xor_0/inv_0/op gnd 0.32fF
C446 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op 0.06fF
C447 gnd ffipg_1/ffi_1/nand_0/w_0_0# 0.10fF
C448 nor_4/b inv_9/in 0.16fF
C449 ffipg_2/ffi_0/inv_1/w_0_6# ffipg_2/ffi_0/inv_1/op 0.04fF
C450 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/ffi_1/q 0.06fF
C451 inv_1/op nor_1/w_0_0# 0.03fF
C452 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C453 cla_2/g1 gnd 0.65fF
C454 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C455 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_3/b 0.00fF
C456 gnd ffipg_0/ffi_1/nand_7/a 0.37fF
C457 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C458 ffipg_1/ffi_0/inv_1/w_0_6# clk 0.06fF
C459 cla_1/inv_0/op cla_0/n 0.06fF
C460 ffi_0/inv_1/op ffi_0/inv_1/w_0_6# 0.04fF
C461 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C462 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_7/a 0.04fF
C463 gnd ffipg_3/ffi_0/nand_0/a_13_n26# 0.01fF
C464 sumffo_0/sbar gnd 0.62fF
C465 nand_2/b cla_0/nand_0/w_0_0# 0.05fF
C466 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C467 sumffo_2/xor_0/inv_1/op ffi_0/q 0.04fF
C468 x3in ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C469 gnd ffipg_0/ffi_0/nand_3/a 0.33fF
C470 gnd inv_9/in 0.33fF
C471 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_1/a 0.04fF
C472 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C473 cla_0/inv_0/in cla_1/p0 0.02fF
C474 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C475 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_0/q 0.06fF
C476 gnd ffipg_0/ffi_0/nand_3/b 0.74fF
C477 gnd sumffo_1/ffo_0/inv_0/op 0.27fF
C478 inv_5/in inv_5/w_0_6# 0.10fF
C479 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C480 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C481 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/b 0.31fF
C482 ffipg_0/k ffipg_0/ffi_0/q 0.07fF
C483 gnd ffipg_2/ffi_1/nand_1/b 0.57fF
C484 gnd ffipg_1/ffi_1/inv_1/op 1.85fF
C485 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# 0.04fF
C486 sumffo_1/ffo_0/nand_1/w_0_0# gnd 0.10fF
C487 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C488 cla_2/p0 gnd 1.06fF
C489 cla_1/l cla_1/nor_0/w_0_0# 0.05fF
C490 inv_0/in nor_0/a 0.02fF
C491 gnd ffipg_0/ffi_1/nand_1/w_0_0# 0.10fF
C492 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C493 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q 0.32fF
C494 gnd ffipg_1/ffi_1/nand_0/a_13_n26# 0.01fF
C495 gnd ffipg_1/ffi_0/nand_1/b 0.57fF
C496 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# 0.04fF
C497 ffi_0/nand_5/w_0_0# ffi_0/nand_1/b 0.06fF
C498 gnd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C499 sumffo_1/ffo_0/nand_6/a clk 0.13fF
C500 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C501 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C502 gnd sumffo_2/ffo_0/nand_2/w_0_0# 0.10fF
C503 gnd cla_0/g0 1.11fF
C504 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/a 0.06fF
C505 ffipg_0/ffi_1/inv_0/op x1in 0.04fF
C506 ffipg_3/ffi_1/inv_0/op ffipg_3/ffi_1/inv_0/w_0_6# 0.03fF
C507 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/qbar 0.00fF
C508 gnd ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C509 sumffo_1/ffo_0/nand_4/w_0_0# clk 0.06fF
C510 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a 0.31fF
C511 gnd ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C512 ffipg_3/ffi_1/q ffipg_3/ffi_0/q 0.73fF
C513 ffi_0/inv_0/op ffi_0/inv_0/w_0_6# 0.03fF
C514 ffipg_1/ffi_0/nand_7/w_0_0# ffipg_1/ffi_0/nand_7/a 0.06fF
C515 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_3/b 0.33fF
C516 cla_1/p0 ffipg_1/ffi_0/q 0.03fF
C517 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# 0.04fF
C518 cla_2/p0 ffipg_2/k 0.05fF
C519 sumffo_0/xor_0/inv_1/op ffi_0/q 0.22fF
C520 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C521 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a 0.31fF
C522 gnd cla_1/inv_0/w_0_6# 0.06fF
C523 ffipg_1/pggen_0/nand_0/w_0_0# ffipg_1/ffi_1/q 0.06fF
C524 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C525 ffipg_3/ffi_1/nand_2/w_0_0# ffipg_3/ffi_1/nand_3/a 0.04fF
C526 sumffo_0/ffo_0/nand_1/b clk 0.45fF
C527 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C528 inv_3/w_0_6# inv_3/in 0.10fF
C529 gnd ffipg_3/ffi_0/nand_7/a 0.37fF
C530 ffipg_0/ffi_1/inv_0/w_0_6# x1in 0.06fF
C531 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C532 ffipg_0/ffi_1/inv_1/w_0_6# clk 0.06fF
C533 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a 0.00fF
C534 gnd z3o 0.80fF
C535 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C536 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# 0.04fF
C537 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C538 gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C539 gnd ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C540 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k 0.06fF
C541 sumffo_0/ffo_0/d clk 0.25fF
C542 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/inv_1/w_0_6# 0.04fF
C543 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C544 gnd ffo_0/nand_3/w_0_0# 0.11fF
C545 sumffo_2/sbar z3o 0.32fF
C546 gnd ffipg_3/ffi_1/nand_3/b 0.74fF
C547 gnd ffipg_2/ffi_1/nand_7/w_0_0# 0.10fF
C548 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_3/b 0.00fF
C549 gnd ffipg_3/ffi_1/nand_6/w_0_0# 0.10fF
C550 ffipg_0/ffi_0/nand_1/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C551 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C552 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C553 gnd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C554 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/inv_0/op 0.06fF
C555 sumffo_2/xor_0/inv_0/w_0_6# inv_1/op 0.06fF
C556 gnd ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C557 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C558 gnd sumffo_1/ffo_0/nand_3/a 0.48fF
C559 nor_0/w_0_0# cla_0/g0 0.06fF
C560 ffi_0/nand_3/b ffi_0/nand_3/a 0.31fF
C561 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_3/b 0.06fF
C562 ffipg_1/ffi_0/q ffipg_1/ffi_1/q 0.73fF
C563 sumffo_3/ffo_0/nand_4/w_0_0# gnd 0.10fF
C564 sumffo_0/ffo_0/inv_0/op gnd 0.27fF
C565 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# 0.16fF
C566 ffipg_2/ffi_1/inv_1/op clk 0.07fF
C567 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C568 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a 0.13fF
C569 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a 0.31fF
C570 gnd ffipg_1/ffi_1/qbar 0.67fF
C571 gnd ffipg_2/ffi_1/nand_6/a 0.37fF
C572 gnd ffipg_0/ffi_0/q 3.00fF
C573 gnd cla_1/inv_0/op 0.27fF
C574 gnd ffipg_3/ffi_1/inv_1/op 1.85fF
C575 ffi_0/nand_6/a nor_0/b 0.00fF
C576 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a 0.00fF
C577 sumffo_1/ffo_0/nand_1/a gnd 0.44fF
C578 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C579 ffi_0/nand_1/a ffi_0/nand_0/w_0_0# 0.04fF
C580 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/nand_1/b 0.06fF
C581 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/q 0.04fF
C582 sumffo_2/ffo_0/inv_1/w_0_6# gnd 0.07fF
C583 gnd ffipg_1/ffi_0/inv_0/op 0.27fF
C584 ffo_0/nand_1/a ffo_0/nand_0/b 0.13fF
C585 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C586 gnd ffo_0/nand_0/b 0.58fF
C587 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a 0.00fF
C588 z3o sumffo_2/ffo_0/nand_7/a 0.00fF
C589 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q 0.32fF
C590 ffipg_0/k ffipg_0/ffi_1/q 0.46fF
C591 ffipg_2/k ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C592 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/qbar 0.31fF
C593 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# 0.04fF
C594 sumffo_2/ffo_0/d gnd 0.41fF
C595 sumffo_0/sbar z1o 0.32fF
C596 ffi_0/nand_1/w_0_0# ffi_0/nand_1/a 0.06fF
C597 gnd ffipg_0/ffi_1/nand_3/a 0.33fF
C598 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_6/a 0.04fF
C599 ffo_0/nand_2/w_0_0# ffo_0/d 0.06fF
C600 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_1/b 0.04fF
C601 gnd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C602 ffipg_0/k nor_0/b 0.06fF
C603 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C604 cla_0/inv_0/in gnd 0.34fF
C605 sumffo_3/ffo_0/nand_7/a sumffo_3/sbar 0.31fF
C606 gnd inv_1/op 0.58fF
C607 ffipg_2/ffi_1/nand_4/w_0_0# ffipg_2/ffi_1/nand_6/a 0.04fF
C608 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C609 sumffo_3/ffo_0/nand_0/b clk 0.04fF
C610 sumffo_2/ffo_0/nand_6/a clk 0.13fF
C611 ffipg_0/ffi_1/inv_0/op ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C612 ffipg_3/ffi_1/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C613 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a 0.00fF
C614 gnd ffo_0/nand_5/w_0_0# 0.10fF
C615 ffipg_1/ffi_0/nand_0/w_0_0# clk 0.06fF
C616 ffipg_0/ffi_0/inv_1/op clk 0.07fF
C617 nand_2/b cla_0/inv_0/op 0.09fF
C618 gnd ffipg_0/ffi_1/nand_2/w_0_0# 0.10fF
C619 clk ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C620 sumffo_1/ffo_0/inv_1/w_0_6# clk 0.06fF
C621 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_1/inv_1/op 0.75fF
C622 ffipg_0/pggen_0/xor_0/inv_0/op gnd 0.32fF
C623 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/op 0.04fF
C624 ffipg_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C625 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C626 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C627 gnd sumffo_3/ffo_0/nand_6/a 0.33fF
C628 cla_0/l inv_2/w_0_6# 0.06fF
C629 y1in ffipg_0/ffi_0/inv_1/op 0.01fF
C630 nand_2/b inv_3/w_0_6# 0.06fF
C631 ffipg_3/ffi_1/nand_7/w_0_0# ffipg_3/ffi_1/nand_7/a 0.06fF
C632 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/inv_1/op 0.06fF
C633 gnd ffipg_1/ffi_0/inv_1/op 1.85fF
C634 gnd ffipg_0/ffi_0/nand_6/w_0_0# 0.10fF
C635 sumffo_1/xor_0/inv_0/op ffi_0/q 0.06fF
C636 ffo_0/nand_2/a_13_n26# gnd 0.01fF
C637 ffipg_3/ffi_0/nand_2/w_0_0# ffipg_3/ffi_0/nand_3/a 0.04fF
C638 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C639 cla_2/g1 cla_2/inv_0/in 0.04fF
C640 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# 0.04fF
C641 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/w_0_0# 0.06fF
C642 ffipg_2/k inv_1/op 0.09fF
C643 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C644 gnd ffipg_1/ffi_0/q 3.00fF
C645 gnd ffi_0/nand_3/a 0.33fF
C646 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a 0.31fF
C647 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C648 gnd ffipg_1/ffi_0/nand_0/a_13_n26# 0.01fF
C649 ffipg_1/ffi_0/nand_6/w_0_0# ffipg_1/ffi_0/nand_6/a 0.06fF
C650 ffipg_0/ffi_1/nand_1/a clk 0.13fF
C651 ffipg_0/ffi_1/nand_1/w_0_0# ffipg_0/ffi_1/nand_3/b 0.04fF
C652 gnd ffo_0/nand_4/w_0_0# 0.10fF
C653 cla_1/l cla_1/p0 0.16fF
C654 cla_0/l cla_1/n 0.13fF
C655 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C656 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C657 ffipg_1/ffi_1/nand_7/w_0_0# gnd 0.10fF
C658 gnd sumffo_3/ffo_0/nand_1/a 0.33fF
C659 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_3/b 0.00fF
C660 ffipg_1/ffi_0/nand_5/w_0_0# ffipg_1/ffi_0/inv_1/op 0.06fF
C661 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C662 ffipg_0/ffi_1/inv_0/op ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C663 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b 0.32fF
C664 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C665 clk ffipg_3/ffi_1/nand_1/a 0.13fF
C666 gnd ffipg_3/ffi_1/nand_3/w_0_0# 0.11fF
C667 ffi_0/nand_1/w_0_0# ffi_0/nand_1/b 0.06fF
C668 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a 0.13fF
C669 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C670 gnd ffipg_0/ffi_1/q 2.24fF
C671 ffipg_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C672 nor_4/b nor_3/w_0_0# 0.03fF
C673 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_3/a 0.04fF
C674 cla_1/l cla_0/n 0.07fF
C675 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C676 gnd ffipg_2/ffi_1/nand_2/w_0_0# 0.10fF
C677 gnd ffo_0/inv_0/op 0.37fF
C678 z3o sumffo_2/ffo_0/nand_7/w_0_0# 0.04fF
C679 cla_0/g0 ffi_0/q 0.08fF
C680 cla_2/l nor_3/b 0.10fF
C681 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a 0.31fF
C682 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# 0.04fF
C683 ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C684 nor_0/b ffi_0/nand_7/w_0_0# 0.06fF
C685 gnd nor_0/b 0.74fF
C686 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C687 gnd sumffo_0/xor_0/a_10_10# 0.93fF
C688 ffipg_2/ffi_0/nand_0/w_0_0# ffipg_2/ffi_0/inv_0/op 0.06fF
C689 ffipg_2/ffi_1/nand_2/w_0_0# ffipg_2/ffi_1/nand_3/a 0.04fF
C690 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C691 ffipg_0/ffi_0/inv_0/op clk 0.32fF
C692 sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# 0.02fF
C693 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C694 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_0/op 0.08fF
C695 gnd nor_3/w_0_0# 0.15fF
C696 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C697 ffipg_0/ffi_1/nand_4/w_0_0# ffipg_0/ffi_1/nand_3/b 0.06fF
C698 ffipg_0/ffi_1/inv_1/op clk 0.07fF
C699 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_3/b 0.31fF
C700 ffo_0/nand_1/b clk 0.45fF
C701 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/qbar 0.04fF
C702 clk ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C703 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C704 ffipg_3/ffi_1/q ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C705 y1in ffipg_0/ffi_0/inv_0/op 0.04fF
C706 y1in clk 0.68fF
C707 gnd ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C708 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C709 sumffo_0/ffo_0/nand_0/b gnd 0.58fF
C710 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_3/b 0.04fF
C711 gnd ffipg_3/ffi_1/nand_1/b 0.57fF
C712 cla_2/n nor_3/b 0.41fF
C713 gnd sumffo_0/xor_0/inv_0/op 0.32fF
C714 gnd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C715 inv_5/w_0_6# cla_0/n 0.06fF
C716 ffo_0/nand_6/w_0_0# ffo_0/nand_6/a 0.06fF
C717 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_1/b 0.45fF
C718 gnd ffipg_1/ffi_1/nand_4/w_0_0# 0.10fF
C719 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/b 0.31fF
C720 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a 0.31fF
C721 ffipg_3/k ffipg_3/ffi_0/q 0.07fF
C722 cla_2/p1 ffipg_3/ffi_0/q 0.03fF
C723 gnd sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C724 gnd sumffo_2/xor_0/w_n3_4# 0.12fF
C725 y3in clk 0.68fF
C726 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a 0.13fF
C727 sumffo_0/xor_0/w_n3_4# gnd 0.12fF
C728 cla_2/g1 cla_2/n 0.13fF
C729 gnd ffipg_2/ffi_0/q 3.00fF
C730 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_1/b 0.45fF
C731 gnd ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C732 ffo_0/d inv_9/in 0.04fF
C733 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C734 cla_2/p0 cla_2/l 0.16fF
C735 nand_2/b cla_0/g0 0.13fF
C736 sumffo_1/xor_0/a_38_n43# ffi_0/q 0.01fF
C737 ffi_0/nand_3/w_0_0# ffi_0/nand_1/b 0.04fF
C738 ffo_0/nand_7/a ffo_0/nand_7/w_0_0# 0.06fF
C739 sumffo_1/ffo_0/nand_5/w_0_0# clk 0.06fF
C740 sumffo_0/ffo_0/nand_4/w_0_0# clk 0.06fF
C741 gnd ffi_0/nand_5/w_0_0# 0.10fF
C742 gnd cla_2/inv_0/w_0_6# 0.06fF
C743 ffipg_1/ffi_1/nand_2/w_0_0# clk 0.06fF
C744 y2in ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C745 inv_6/in nor_4/b 0.04fF
C746 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b 0.13fF
C747 gnd ffipg_3/ffi_0/nand_2/w_0_0# 0.10fF
C748 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/inv_1/op 0.13fF
C749 sumffo_3/ffo_0/inv_0/op gnd 0.52fF
C750 ffipg_1/ffi_0/nand_4/w_0_0# ffipg_1/ffi_0/nand_3/b 0.06fF
C751 gnd ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C752 cla_2/p0 ffipg_2/ffi_1/q 0.22fF
C753 gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C754 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C755 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C756 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/inv_0/w_0_6# 0.03fF
C757 nor_0/w_0_0# nor_0/b 0.06fF
C758 ffo_0/qbar couto 0.32fF
C759 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C760 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/inv_1/w_0_6# 0.04fF
C761 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/inv_1/op 0.33fF
C762 ffipg_2/k ffipg_2/ffi_0/q 0.07fF
C763 sumffo_3/ffo_0/nand_6/w_0_0# gnd 0.10fF
C764 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/nand_7/a 0.04fF
C765 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C766 inv_6/in gnd 0.33fF
C767 gnd sumffo_3/ffo_0/nand_2/w_0_0# 0.10fF
C768 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C769 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_3/b 0.31fF
C770 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C771 sumffo_2/ffo_0/inv_0/w_0_6# gnd 0.07fF
C772 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/op 0.04fF
C773 gnd ffipg_0/ffi_0/nand_6/a 0.37fF
C774 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_3/a 0.06fF
C775 inv_1/in nor_1/b 0.16fF
C776 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C777 ffi_0/inv_1/op ffi_0/nand_1/b 0.45fF
C778 cla_0/l cla_1/p0 0.09fF
C779 gnd ffipg_2/ffi_0/nand_0/a_13_n26# 0.01fF
C780 gnd cla_1/nand_0/a_13_n26# 0.01fF
C781 gnd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C782 ffi_0/nand_2/w_0_0# clk 0.06fF
C783 gnd ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C784 y4in ffipg_3/ffi_0/inv_1/op 0.01fF
C785 sumffo_2/ffo_0/d ffi_0/q 0.27fF
C786 clk ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C787 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C788 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C789 cla_0/l inv_7/w_0_6# 0.06fF
C790 gnd ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C791 sumffo_3/xor_0/inv_0/w_0_6# gnd 0.09fF
C792 cla_1/l gnd 0.40fF
C793 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C794 ffipg_3/k cla_0/l 0.10fF
C795 sumffo_1/ffo_0/nand_1/b clk 0.45fF
C796 sumffo_2/ffo_0/inv_0/w_0_6# sumffo_2/ffo_0/inv_0/op 0.03fF
C797 cla_0/l cla_2/p1 0.30fF
C798 cla_1/nand_0/w_0_0# cla_0/l 0.06fF
C799 cla_0/l cla_0/n 0.25fF
C800 cla_0/g0 nor_0/a 0.68fF
C801 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a 0.13fF
C802 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C803 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/nand_7/a 0.06fF
C804 ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C805 gnd ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C806 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar 0.32fF
C807 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C808 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# 0.04fF
C809 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C810 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a 0.00fF
C811 ffipg_1/ffi_1/nand_0/w_0_0# clk 0.06fF
C812 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_0/q 0.12fF
C813 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.35fF
C814 gnd ffipg_1/ffi_1/nand_1/a 0.44fF
C815 ffipg_0/ffi_0/nand_2/w_0_0# ffipg_0/ffi_0/nand_3/a 0.04fF
C816 sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d 0.52fF
C817 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C818 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# 0.04fF
C819 gnd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C820 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_1/w_0_6# 0.03fF
C821 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# 0.04fF
C822 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C823 gnd ffipg_0/ffi_1/nand_3/w_0_0# 0.11fF
C824 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a 0.00fF
C825 gnd inv_5/w_0_6# 0.42fF
C826 ffi_0/nand_1/w_0_0# ffi_0/nand_3/b 0.04fF
C827 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/q 0.31fF
C828 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C829 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C830 gnd ffipg_3/ffi_0/qbar 0.67fF
C831 gnd ffipg_2/ffi_1/nand_7/a 0.37fF
C832 ffipg_1/ffi_1/inv_0/op x2in 0.04fF
C833 gnd cla_1/inv_0/in 0.34fF
C834 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/qbar 0.04fF
C835 gnd ffipg_3/ffi_1/nand_6/a 0.37fF
C836 gnd ffipg_3/ffi_0/q 3.00fF
C837 ffipg_0/ffi_0/nand_3/a clk 0.13fF
C838 ffipg_2/ffi_1/nand_0/w_0_0# ffipg_2/ffi_1/inv_0/op 0.06fF
C839 x2in ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C840 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a 0.31fF
C841 gnd ffi_0/inv_1/w_0_6# 0.06fF
C842 ffo_0/d ffo_0/nand_0/b 0.40fF
C843 ffipg_0/ffi_0/inv_1/w_0_6# ffipg_0/ffi_0/inv_1/op 0.04fF
C844 ffi_0/nand_1/a ffi_0/nand_1/b 0.31fF
C845 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C846 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/qbar 0.00fF
C847 ffipg_1/ffi_1/inv_1/op clk 0.07fF
C848 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C849 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a 0.31fF
C850 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/a 0.06fF
C851 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_3/a 0.04fF
C852 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_1/a 0.06fF
C853 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/qbar 0.31fF
C854 ffi_0/inv_0/op cinin 0.04fF
C855 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C856 gnd ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C857 sumffo_2/ffo_0/nand_1/b gnd 0.57fF
C858 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/inv_1/w_0_6# 0.04fF
C859 nor_4/a inv_8/in 0.04fF
C860 ffipg_1/ffi_0/inv_0/op ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C861 gnd cla_2/nor_0/w_0_0# 0.31fF
C862 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q 0.22fF
C863 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op 0.13fF
C864 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C865 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_1/b 0.31fF
C866 gnd ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C867 nor_0/a ffipg_0/ffi_0/q 0.03fF
C868 nor_4/a inv_8/w_0_6# 0.03fF
C869 inv_7/op inv_7/w_0_6# 0.03fF
C870 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# 0.04fF
C871 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C872 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_3/b 0.00fF
C873 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/ffi_0/q 0.23fF
C874 ffi_0/nand_6/w_0_0# ffi_0/nand_6/a 0.06fF
C875 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C876 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/q 0.31fF
C877 gnd x1in 0.22fF
C878 nor_0/b ffi_0/q 0.32fF
C879 sumffo_0/xor_0/a_10_10# ffi_0/q 0.12fF
C880 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C881 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a 0.00fF
C882 gnd sumffo_0/ffo_0/nand_7/a 0.33fF
C883 ffi_0/nand_3/b ffi_0/nand_3/w_0_0# 0.06fF
C884 gnd ffi_0/nand_0/w_0_0# 0.10fF
C885 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/nand_6/a 0.06fF
C886 gnd y2in 0.22fF
C887 gnd ffipg_0/ffi_0/qbar 0.67fF
C888 inv_7/op inv_8/w_0_6# 0.06fF
C889 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C890 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/a 0.06fF
C891 ffi_0/inv_1/op ffi_0/nand_6/a 0.13fF
C892 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C893 ffo_0/nand_3/a ffo_0/nand_3/w_0_0# 0.06fF
C894 inv_2/in inv_2/w_0_6# 0.10fF
C895 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_3/b 0.00fF
C896 ffipg_2/ffi_0/nand_1/a gnd 0.44fF
C897 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C898 ffi_0/inv_0/op gnd 0.27fF
C899 gnd ffipg_0/ffi_1/nand_7/w_0_0# 0.10fF
C900 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C901 sumffo_0/xor_0/inv_0/op ffi_0/q 0.20fF
C902 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_7/a 0.04fF
C903 gnd ffipg_1/ffi_0/nand_3/b 0.74fF
C904 inv_0/in nor_0/b 0.16fF
C905 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C906 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_1/op 0.52fF
C907 ffipg_0/ffi_1/nand_4/w_0_0# ffipg_0/ffi_1/inv_1/op 0.06fF
C908 gnd x4in 0.22fF
C909 ffi_0/nand_1/w_0_0# gnd 0.10fF
C910 nor_4/a nor_4/w_0_0# 0.07fF
C911 gnd cla_0/l 3.05fF
C912 x3in ffipg_2/ffi_1/inv_0/op 0.04fF
C913 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C914 sumffo_2/xor_0/w_n3_4# ffi_0/q 0.00fF
C915 ffo_0/nand_1/b ffo_0/nand_3/w_0_0# 0.04fF
C916 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C917 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C918 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C919 sumffo_2/ffo_0/nand_3/a gnd 0.33fF
C920 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C921 sumffo_0/xor_0/w_n3_4# ffi_0/q 0.06fF
C922 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op 0.06fF
C923 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C924 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C925 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C926 ffipg_2/ffi_1/nand_5/w_0_0# ffipg_2/ffi_1/nand_7/a 0.04fF
C927 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/b 0.31fF
C928 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C929 ffipg_0/ffi_0/inv_1/w_0_6# clk 0.06fF
C930 sumffo_3/ffo_0/nand_4/w_0_0# clk 0.06fF
C931 gnd cla_0/nor_1/w_0_0# 0.31fF
C932 sumffo_0/xor_0/w_n3_4# sumffo_0/ffo_0/d 0.02fF
C933 ffi_0/nand_3/b ffi_0/inv_1/op 0.33fF
C934 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C935 inv_5/in cla_0/n 0.13fF
C936 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C937 clk ffipg_3/ffi_1/inv_1/op 0.07fF
C938 ffo_0/d ffo_0/inv_0/op 0.04fF
C939 ffo_0/nand_1/w_0_0# ffo_0/nand_1/a 0.06fF
C940 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b 0.13fF
C941 ffipg_2/k cla_0/l 0.10fF
C942 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C943 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C944 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C945 ffo_0/nand_3/a ffo_0/nand_0/b 0.13fF
C946 gnd ffo_0/nand_1/w_0_0# 0.10fF
C947 sumffo_3/xor_0/a_10_10# sumffo_3/ffo_0/d 0.45fF
C948 sumffo_1/xor_0/inv_1/w_0_6# gnd 0.06fF
C949 gnd cla_0/inv_0/w_0_6# 0.06fF
C950 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_1/b 0.04fF
C951 sumffo_2/ffo_0/inv_1/w_0_6# clk 0.06fF
C952 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C953 ffipg_1/ffi_0/inv_0/op clk 0.32fF
C954 ffipg_3/ffi_0/inv_0/op y4in 0.04fF
C955 ffo_0/nand_0/b clk 0.04fF
C956 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/w_0_0# 0.06fF
C957 gnd ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C958 gnd ffipg_1/ffi_1/nand_3/b 0.74fF
C959 nor_4/b nor_4/a 0.42fF
C960 ffo_0/nand_3/b ffo_0/nand_1/a 0.00fF
C961 sumffo_1/sbar z2o 0.32fF
C962 ffipg_2/ffi_0/nand_2/w_0_0# ffipg_2/ffi_0/nand_3/a 0.04fF
C963 gnd ffo_0/nand_3/b 0.74fF
C964 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_1/b 0.45fF
C965 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C966 nor_2/b cla_1/n 0.39fF
C967 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C968 ffipg_3/k ffipg_3/ffi_1/q 0.46fF
C969 cla_2/p1 ffipg_3/ffi_1/q 0.22fF
C970 cinin ffi_0/inv_0/w_0_6# 0.06fF
C971 cla_1/nor_0/w_0_0# cla_1/p0 0.06fF
C972 sumffo_2/ffo_0/d clk 0.25fF
C973 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# 0.04fF
C974 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/d 0.40fF
C975 sumffo_0/ffo_0/inv_0/w_0_6# gnd 0.06fF
C976 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_1/b 0.06fF
C977 ffipg_1/k cla_1/p0 0.05fF
C978 ffipg_0/ffi_1/nand_3/a clk 0.13fF
C979 gnd sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C980 gnd ffipg_1/ffi_1/nand_7/a 0.37fF
C981 gnd ffipg_1/ffi_0/nand_3/a 0.33fF
C982 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C983 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C984 cinin ffi_0/inv_1/op 0.01fF
C985 gnd ffi_0/nand_3/w_0_0# 0.11fF
C986 cla_2/n nor_3/w_0_0# 0.06fF
C987 inv_1/in inv_1/op 0.04fF
C988 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C989 gnd cla_1/nor_1/w_0_0# 0.31fF
C990 cla_0/l inv_7/in 0.13fF
C991 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/ffi_1/q 0.06fF
C992 sumffo_3/ffo_0/nand_7/a gnd 0.33fF
C993 sumffo_0/ffo_0/nand_5/w_0_0# gnd 0.10fF
C994 nor_0/b ffi_0/nand_7/a 0.31fF
C995 gnd nor_4/a 0.40fF
C996 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C997 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/a 0.31fF
C998 nor_0/a ffipg_0/ffi_1/q 0.22fF
C999 gnd ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1000 ffo_0/nand_5/w_0_0# clk 0.06fF
C1001 gnd sumffo_0/ffo_0/nand_7/w_0_0# 0.10fF
C1002 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C1003 sumffo_3/ffo_0/nand_7/a z4o 0.00fF
C1004 ffipg_2/ffi_1/nand_0/w_0_0# gnd 0.10fF
C1005 gnd ffipg_2/ffi_0/inv_1/op 1.85fF
C1006 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_0/q 0.20fF
C1007 gnd inv_0/op 0.27fF
C1008 ffipg_0/ffi_1/nand_2/w_0_0# clk 0.06fF
C1009 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C1010 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_3/b 0.06fF
C1011 ffipg_1/ffi_1/inv_0/op ffipg_1/ffi_1/inv_0/w_0_6# 0.03fF
C1012 x4in ffipg_3/ffi_1/inv_0/op 0.04fF
C1013 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C1014 sumffo_3/ffo_0/nand_6/a clk 0.13fF
C1015 gnd sumffo_1/xor_0/w_n3_4# 0.12fF
C1016 gnd ffipg_0/ffi_1/nand_0/w_0_0# 0.10fF
C1017 gnd ffi_0/nand_6/w_0_0# 0.10fF
C1018 nor_0/a nor_0/b 0.32fF
C1019 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# 0.16fF
C1020 gnd inv_7/op 0.27fF
C1021 ffipg_2/ffi_1/q ffipg_2/ffi_0/q 0.73fF
C1022 ffipg_1/ffi_0/inv_1/op clk 0.07fF
C1023 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C1024 ffi_0/nand_1/a ffi_0/nand_3/b 0.00fF
C1025 gnd ffi_0/inv_0/w_0_6# 0.06fF
C1026 gnd ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C1027 gnd ffipg_2/ffi_0/nand_3/a 0.33fF
C1028 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C1029 gnd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C1030 ffipg_1/ffi_0/nand_7/w_0_0# ffipg_1/ffi_0/q 0.04fF
C1031 gnd sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C1032 gnd ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C1033 ffipg_2/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C1034 gnd ffo_0/nand_7/a 0.33fF
C1035 ffo_0/nand_6/w_0_0# gnd 0.10fF
C1036 ffi_0/nand_3/a clk 0.13fF
C1037 ffo_0/inv_0/op ffo_0/inv_0/w_0_6# 0.03fF
C1038 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C1039 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q 0.22fF
C1040 gnd sumffo_3/ffo_0/d 0.41fF
C1041 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C1042 ffipg_1/k ffipg_1/ffi_1/q 0.46fF
C1043 gnd ffipg_0/ffi_1/inv_0/op 0.27fF
C1044 sumffo_3/xor_0/inv_1/w_0_6# gnd 0.06fF
C1045 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C1046 ffi_0/nand_5/w_0_0# ffi_0/nand_7/a 0.04fF
C1047 gnd ffi_0/inv_1/op 1.89fF
C1048 z1o sumffo_0/ffo_0/nand_7/a 0.00fF
C1049 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/d 0.06fF
C1050 nand_2/b cla_1/l 0.31fF
C1051 ffo_0/nand_4/w_0_0# clk 0.06fF
C1052 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/inv_1/w_0_6# 0.04fF
C1053 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1054 cla_0/inv_0/in cla_0/inv_0/op 0.04fF
C1055 gnd y4in 0.22fF
C1056 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C1057 gnd z2o 0.80fF
C1058 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/ffi_0/q 0.06fF
C1059 gnd sumffo_3/sbar 0.62fF
C1060 gnd sumffo_0/ffo_0/nand_1/a 0.44fF
C1061 ffipg_2/ffi_0/inv_0/w_0_6# ffipg_2/ffi_0/inv_0/op 0.03fF
C1062 sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d 0.06fF
C1063 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# 0.16fF
C1064 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1065 ffipg_2/k sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C1066 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C1067 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C1068 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C1069 inv_6/in cla_2/n 0.02fF
C1070 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a 0.31fF
C1071 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C1072 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C1073 gnd x2in 0.22fF
C1074 sumffo_3/sbar z4o 0.32fF
C1075 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar 0.32fF
C1076 ffipg_0/pggen_0/nand_0/w_0_0# gnd 0.10fF
C1077 gnd ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C1078 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C1079 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C1080 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_1/b 0.04fF
C1081 ffipg_2/ffi_1/nand_2/w_0_0# clk 0.06fF
C1082 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_1/b 0.31fF
C1083 ffipg_2/ffi_1/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C1084 gnd sumffo_2/ffo_0/nand_3/w_0_0# 0.11fF
C1085 inv_5/in gnd 0.49fF
C1086 inv_0/op nor_0/w_0_0# 0.10fF
C1087 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_3/b 0.04fF
C1088 ffipg_2/ffi_1/nand_1/a gnd 0.44fF
C1089 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C1090 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C1091 gnd x3in 0.22fF
C1092 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a 0.13fF
C1093 ffo_0/inv_1/w_0_6# gnd 0.06fF
C1094 ffipg_3/ffi_1/q ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1095 inv_7/op inv_7/in 0.04fF
C1096 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_1/b 0.31fF
C1097 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C1098 cla_2/l inv_5/w_0_6# 0.08fF
C1099 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C1100 gnd ffipg_3/ffi_1/q 2.24fF
C1101 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_0/op 0.08fF
C1102 gnd sumffo_0/ffo_0/nand_1/w_0_0# 0.10fF
C1103 ffi_0/nand_3/b ffi_0/nand_1/b 0.32fF
C1104 ffipg_2/ffi_0/nand_4/w_0_0# gnd 0.10fF
C1105 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_1/w_0_0# 0.06fF
C1106 sumffo_0/ffo_0/nand_0/b clk 0.04fF
C1107 ffo_0/nand_0/w_0_0# ffo_0/nand_1/a 0.04fF
C1108 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a 0.13fF
C1109 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op 0.13fF
C1110 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a 0.31fF
C1111 gnd ffo_0/nand_0/w_0_0# 0.10fF
C1112 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1113 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1114 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C1115 gnd ffi_0/nand_1/a 0.44fF
C1116 sumffo_3/xor_0/inv_1/op ffipg_3/k 0.22fF
C1117 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1118 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C1119 cla_0/l cla_2/inv_0/in 0.16fF
C1120 gnd ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C1121 gnd cla_1/nor_0/w_0_0# 0.31fF
C1122 ffi_0/nand_2/w_0_0# ffi_0/nand_3/a 0.04fF
C1123 ffipg_1/ffi_0/nand_6/w_0_0# ffipg_1/ffi_0/q 0.06fF
C1124 ffipg_1/k gnd 0.70fF
C1125 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_1/b 0.04fF
C1126 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1127 cla_0/g0 ffipg_0/ffi_0/q 0.13fF
C1128 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a 0.00fF
C1129 cla_0/l ffi_0/q 0.33fF
C1130 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.35fF
C1131 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_7/w_0_0# 0.06fF
C1132 gnd sumffo_1/ffo_0/d 0.41fF
C1133 gnd ffo_0/nand_6/a 0.33fF
C1134 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/ffi_0/q 0.06fF
C1135 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C1136 clk ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1137 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C1138 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C1139 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# 0.04fF
C1140 z1o sumffo_0/ffo_0/nand_7/w_0_0# 0.04fF
C1141 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a 0.00fF
C1142 gnd inv_2/w_0_6# 0.17fF
C1143 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/qbar 0.00fF
C1144 gnd ffipg_0/ffi_0/nand_0/w_0_0# 0.10fF
C1145 ffipg_2/ffi_0/nand_0/w_0_0# clk 0.06fF
C1146 sumffo_3/xor_0/inv_1/op inv_4/op 0.06fF
C1147 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C1148 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_1/q 0.06fF
C1149 gnd ffo_0/nand_7/w_0_0# 0.10fF
C1150 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C1151 gnd ffipg_2/ffi_1/qbar 0.67fF
C1152 nor_1/w_0_0# cla_0/n 0.06fF
C1153 cla_2/nor_1/w_0_0# cla_0/l 0.06fF
C1154 cla_0/inv_0/in cla_0/g0 0.16fF
C1155 sumffo_2/ffo_0/nand_6/w_0_0# gnd 0.10fF
C1156 nand_2/b cla_0/l 0.06fF
C1157 gnd ffipg_0/ffi_0/nand_7/w_0_0# 0.10fF
C1158 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C1159 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C1160 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_0/q 0.20fF
C1161 gnd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C1162 sumffo_1/xor_0/a_10_10# sumffo_1/ffo_0/d 0.45fF
C1163 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C1164 gnd cla_1/n 0.51fF
C1165 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/inv_1/op 0.33fF
C1166 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a 0.31fF
C1167 gnd sumffo_2/ffo_0/nand_0/w_0_0# 0.10fF
C1168 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_0/inv_1/op 0.75fF
C1169 gnd ffipg_1/ffi_0/nand_1/a 0.44fF
C1170 ffipg_1/ffi_1/nand_3/a gnd 0.33fF
C1171 gnd ffipg_3/ffi_0/inv_1/op 1.85fF
C1172 ffipg_2/ffi_1/inv_1/w_0_6# clk 0.06fF
C1173 cla_0/l cla_2/l 0.37fF
C1174 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# 0.04fF
C1175 gnd ffi_0/nand_1/b 0.57fF
C1176 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/inv_1/op 0.45fF
C1177 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C1178 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a 0.00fF
C1179 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C1180 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1181 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C1182 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a 0.13fF
C1183 ffipg_3/k cla_2/p1 0.05fF
C1184 ffipg_3/k cla_0/n 0.06fF
C1185 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/nand_6/a 0.04fF
C1186 gnd ffipg_0/ffi_1/nand_1/b 0.57fF
C1187 nor_3/b nor_3/w_0_0# 0.06fF
C1188 sumffo_1/ffo_0/nand_6/w_0_0# z2o 0.06fF
C1189 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C1190 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a 0.13fF
C1191 cla_0/l cla_0/nand_0/w_0_0# 0.06fF
C1192 inv_2/in gnd 0.47fF
C1193 ffipg_1/ffi_1/nand_1/a clk 0.13fF
C1194 cla_1/p0 ffipg_1/ffi_1/q 0.22fF
C1195 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C1196 sumffo_1/xor_0/w_n3_4# ffi_0/q 0.00fF
C1197 inv_8/in inv_8/w_0_6# 0.10fF
C1198 ffi_0/nand_6/w_0_0# ffi_0/q 0.06fF
C1199 inv_7/op ffi_0/q 0.31fF
C1200 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a 0.13fF
C1201 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C1202 sumffo_1/ffo_0/nand_6/a z2o 0.31fF
C1203 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C1204 gnd sumffo_0/ffo_0/nand_6/a 0.33fF
C1205 gnd ffipg_1/ffi_1/inv_0/op 0.27fF
C1206 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# 0.04fF
C1207 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_1/b 0.45fF
C1208 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b 0.32fF
C1209 sumffo_3/xor_0/w_n3_4# sumffo_3/ffo_0/d 0.02fF
C1210 sumffo_1/ffo_0/nand_2/a_13_n26# gnd 0.01fF
C1211 gnd ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C1212 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a 0.13fF
C1213 inv_0/in inv_0/op 0.04fF
C1214 sumffo_3/xor_0/inv_1/op gnd 0.35fF
C1215 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C1216 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/xor_0/inv_0/op 0.03fF
C1217 gnd sumffo_2/ffo_0/nand_3/b 0.74fF
C1218 ffipg_2/ffi_1/nand_1/w_0_0# gnd 0.10fF
C1219 sumffo_3/ffo_0/d ffi_0/q 0.16fF
C1220 clk ffi_0/inv_1/w_0_6# 0.06fF
C1221 inv_4/op ffipg_3/k 0.09fF
C1222 gnd ffipg_3/ffi_0/nand_1/a 0.44fF
C1223 gnd nor_2/b 0.32fF
C1224 sumffo_3/ffo_0/nand_0/w_0_0# gnd 0.10fF
C1225 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# 0.04fF
C1226 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a 0.13fF
C1227 sumffo_3/xor_0/a_10_10# ffipg_3/k 0.12fF
C1228 cla_0/l nor_0/a 0.16fF
C1229 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/w_0_0# 0.04fF
C1230 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/ffi_1/q 0.06fF
C1231 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# 0.04fF
C1232 ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_1/inv_1/op 0.75fF
C1233 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C1234 cla_2/nand_0/w_0_0# gnd 0.18fF
C1235 cla_1/l inv_3/w_0_6# 0.06fF
C1236 ffipg_0/ffi_0/nand_4/w_0_0# gnd 0.10fF
C1237 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_6/a 0.04fF
C1238 gnd sumffo_3/ffo_0/nand_3/a 0.33fF
C1239 sumffo_2/ffo_0/nand_0/b gnd 0.63fF
C1240 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C1241 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# 0.16fF
C1242 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C1243 ffipg_2/ffi_0/inv_1/w_0_6# clk 0.06fF
C1244 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_0/q 0.20fF
C1245 sumffo_2/ffo_0/nand_1/b clk 0.45fF
C1246 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C1247 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1248 nor_2/w_0_0# cla_1/n 0.06fF
C1249 gnd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C1250 ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C1251 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C1252 gnd ffipg_0/ffi_0/nand_1/b 0.57fF
C1253 gnd ffipg_1/ffi_0/nand_4/w_0_0# 0.10fF
C1254 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C1255 inv_6/in nor_3/b 0.16fF
C1256 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C1257 gnd nor_1/w_0_0# 0.15fF
C1258 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C1259 gnd ffipg_2/ffi_1/nand_3/b 0.74fF
C1260 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_3/b 0.00fF
C1261 cla_2/p0 ffipg_2/ffi_0/q 0.03fF
C1262 sumffo_2/xor_0/inv_0/op gnd 0.32fF
C1263 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/b 0.31fF
C1264 gnd ffipg_1/ffi_0/nand_2/w_0_0# 0.10fF
C1265 x1in clk 0.68fF
C1266 gnd ffipg_2/ffi_1/inv_0/op 0.27fF
C1267 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_3/a 0.06fF
C1268 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C1269 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_0/op 0.32fF
C1270 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# 0.04fF
C1271 gnd ffi_0/nand_0/a_13_n26# 0.01fF
C1272 ffi_0/nand_0/w_0_0# clk 0.06fF
C1273 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C1274 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a 0.13fF
C1275 y2in clk 0.68fF
C1276 ffipg_0/ffi_1/inv_1/op x1in 0.01fF
C1277 sumffo_1/ffo_0/nand_0/b gnd 0.62fF
C1278 gnd ffipg_0/ffi_0/nand_3/w_0_0# 0.11fF
C1279 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a 0.31fF
C1280 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/qbar 0.06fF
C1281 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C1282 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_3/b 0.00fF
C1283 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C1284 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1285 ffipg_2/ffi_0/nand_1/a clk 0.13fF
C1286 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C1287 gnd cla_1/p0 1.06fF
C1288 ffi_0/inv_0/op clk 0.32fF
C1289 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C1290 gnd ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C1291 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_7/a 0.04fF
C1292 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C1293 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/ffi_1/q 0.06fF
C1294 gnd ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1295 gnd inv_7/w_0_6# 0.15fF
C1296 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_6/a 0.04fF
C1297 clk x4in 0.68fF
C1298 gnd ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C1299 gnd ffi_0/nand_6/a 0.33fF
C1300 ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C1301 ffipg_2/k sumffo_2/xor_0/inv_0/op 0.20fF
C1302 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C1303 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1304 ffipg_0/ffi_0/q ffipg_0/ffi_1/q 0.73fF
C1305 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C1306 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C1307 gnd ffipg_2/ffi_0/nand_7/a 0.37fF
C1308 ffipg_3/k gnd 0.61fF
C1309 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b 0.13fF
C1310 gnd cla_2/p1 1.00fF
C1311 gnd inv_8/in 0.43fF
C1312 gnd cla_0/n 1.18fF
C1313 ffipg_1/k ffi_0/q 0.06fF
C1314 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b 0.32fF
C1315 gnd ffipg_3/ffi_0/nand_3/a 0.33fF
C1316 ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1317 cla_1/nand_0/w_0_0# gnd 0.10fF
C1318 x3in ffipg_2/ffi_1/inv_1/op 0.01fF
C1319 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/ffi_1/q 0.06fF
C1320 inv_5/in cla_2/l 0.05fF
C1321 sumffo_1/ffo_0/d ffi_0/q 0.27fF
C1322 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/nand_6/a 0.06fF
C1323 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_1/a 0.06fF
C1324 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_0/b 0.40fF
C1325 ffipg_2/k cla_1/p0 0.06fF
C1326 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C1327 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/nand_1/a 0.04fF
C1328 sumffo_1/ffo_0/nand_7/a sumffo_1/sbar 0.31fF
C1329 gnd inv_8/w_0_6# 0.15fF
C1330 nor_2/w_0_0# nor_2/b 0.06fF
C1331 ffo_0/nand_0/b ffo_0/inv_0/op 0.32fF
C1332 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C1333 nor_3/b inv_5/w_0_6# 0.17fF
C1334 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C1335 ffipg_3/ffi_0/nand_4/w_0_0# ffipg_3/ffi_0/inv_1/op 0.06fF
C1336 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C1337 cla_2/p0 cla_1/l 0.02fF
C1338 inv_2/w_0_6# ffi_0/q 0.06fF
C1339 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_0/op 0.32fF
C1340 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_0/q 0.20fF
C1341 nor_4/b nor_4/w_0_0# 0.06fF
C1342 ffipg_0/k gnd 0.68fF
C1343 cla_0/nand_0/a_13_n26# gnd 0.00fF
C1344 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# 0.04fF
C1345 ffo_0/nand_3/b ffo_0/nand_3/a 0.31fF
C1346 gnd ffi_0/nand_3/b 0.74fF
C1347 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/qbar 0.04fF
C1348 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/b 0.31fF
C1349 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C1350 gnd ffipg_1/ffi_1/q 2.24fF
C1351 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# 0.04fF
C1352 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C1353 ffipg_2/k cla_0/n 0.06fF
C1354 gnd ffipg_3/ffi_0/inv_0/op 0.27fF
C1355 ffo_0/nand_3/b clk 0.33fF
C1356 inv_4/op gnd 0.58fF
C1357 z1o sumffo_0/ffo_0/nand_6/a 0.31fF
C1358 gnd sumffo_0/ffo_0/nand_6/w_0_0# 0.10fF
C1359 gnd sumffo_0/ffo_0/nand_3/w_0_0# 0.11fF
C1360 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_1/b 0.45fF
C1361 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C1362 cla_2/g1 ffipg_3/ffi_0/q 0.13fF
C1363 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C1364 sumffo_3/ffo_0/nand_3/b gnd 0.74fF
C1365 gnd sumffo_1/sbar 0.62fF
C1366 sumffo_3/xor_0/a_10_10# gnd 0.93fF
C1367 nand_2/b ffipg_1/k 0.15fF
C1368 ffo_0/nand_3/b ffo_0/nand_1/b 0.32fF
C1369 sumffo_0/ffo_0/inv_1/w_0_6# clk 0.06fF
C1370 cla_0/l cla_0/inv_0/op 0.35fF
C1371 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/inv_1/op 0.33fF
C1372 ffipg_1/ffi_0/nand_3/a clk 0.13fF
C1373 gnd nor_4/w_0_0# 0.15fF
C1374 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C1375 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q 0.27fF
C1376 gnd ffipg_1/ffi_1/nand_5/w_0_0# 0.10fF
C1377 nor_2/b inv_3/in 0.04fF
C1378 inv_7/in inv_7/w_0_6# 0.10fF
C1379 nor_4/a clk 0.03fF
C1380 gnd ffipg_2/ffi_0/inv_0/op 0.27fF
C1381 ffipg_1/ffi_0/qbar gnd 0.67fF
C1382 sumffo_3/xor_0/inv_0/op inv_4/op 0.27fF
C1383 sumffo_0/ffo_0/nand_5/w_0_0# clk 0.06fF
C1384 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1385 ffipg_1/ffi_0/inv_0/op ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C1386 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b 0.32fF
C1387 ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C1388 nand_2/b inv_2/w_0_6# 0.03fF
C1389 gnd ffipg_2/ffi_0/nand_2/w_0_0# 0.10fF
C1390 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a 0.13fF
C1391 ffipg_1/ffi_1/inv_1/w_0_6# clk 0.06fF
C1392 cla_2/p0 cla_1/inv_0/in 0.02fF
C1393 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a 0.31fF
C1394 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b 0.32fF
C1395 ffipg_2/ffi_1/nand_0/w_0_0# clk 0.06fF
C1396 ffipg_2/ffi_0/inv_1/op clk 0.07fF
C1397 sumffo_2/xor_0/inv_0/w_0_6# gnd 0.09fF
C1398 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C1399 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C1400 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar 0.32fF
C1401 gnd cinin 0.22fF
C1402 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C1403 gnd ffipg_0/ffi_0/nand_7/a 0.37fF
C1404 gnd ffipg_1/ffi_1/nand_6/w_0_0# 0.10fF
C1405 ffipg_0/ffi_1/nand_0/w_0_0# clk 0.06fF
C1406 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C1407 sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d 0.52fF
C1408 cla_2/inv_0/op gnd 0.27fF
C1409 cla_0/inv_0/w_0_6# cla_0/inv_0/op 0.03fF
C1410 x4in ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C1411 ffipg_3/ffi_1/nand_2/w_0_0# x4in 0.06fF
C1412 ffo_0/qbar ffo_0/nand_7/a 0.31fF
C1413 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1414 ffo_0/nand_6/w_0_0# ffo_0/qbar 0.04fF
C1415 gnd ffipg_2/ffi_0/nand_1/b 0.57fF
C1416 ffipg_2/ffi_0/nand_3/a clk 0.13fF
C1417 inv_2/in ffi_0/q 0.13fF
C1418 sumffo_3/ffo_0/inv_1/w_0_6# clk 0.06fF
C1419 sumffo_1/ffo_0/nand_7/a gnd 0.33fF
C1420 nor_4/b gnd 0.25fF
C1421 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_3/b 0.04fF
C1422 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a 0.31fF
C1423 ffipg_2/ffi_0/inv_1/op y3in 0.01fF
C1424 sumffo_3/ffo_0/d clk 0.04fF
C1425 gnd ffipg_2/ffi_0/nand_5/w_0_0# 0.10fF
C1426 ffipg_0/ffi_1/inv_0/op clk 0.32fF
C1427 ffo_0/nand_1/b ffo_0/nand_7/a 0.13fF
C1428 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C1429 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C1430 cla_1/inv_0/in cla_1/inv_0/w_0_6# 0.06fF
C1431 clk ffi_0/inv_1/op 0.93fF
C1432 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C1433 sumffo_0/sbar sumffo_0/ffo_0/nand_7/a 0.31fF
C1434 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C1435 gnd sumffo_2/ffo_0/nand_4/w_0_0# 0.10fF
C1436 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/ffi_0/q 0.06fF
C1437 sumffo_3/xor_0/inv_1/op ffi_0/q 0.04fF
C1438 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a 0.31fF
C1439 clk y4in 0.64fF
C1440 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C1441 gnd ffo_0/nand_1/a 0.33fF
C1442 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/d 0.06fF
C1443 sumffo_2/ffo_0/nand_5/w_0_0# gnd 0.10fF
C1444 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a 0.00fF
C1445 gnd ffi_0/nand_7/w_0_0# 0.10fF
C1446 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1447 sumffo_1/ffo_0/nand_3/b gnd 0.74fF
C1448 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C1449 cla_2/g1 cla_0/l 0.26fF
C1450 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C1451 ffipg_1/k nor_0/a 0.06fF
C1452 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C1453 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar 0.32fF
C1454 x2in clk 0.68fF
C1455 ffi_0/nand_4/w_0_0# ffi_0/inv_1/op 0.06fF
C1456 inv_4/op nor_2/w_0_0# 0.03fF
C1457 sumffo_3/ffo_0/inv_0/w_0_6# gnd 0.07fF
C1458 gnd z4o 0.80fF
C1459 gnd sumffo_2/sbar 0.62fF
C1460 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/w_0_0# 0.06fF
C1461 nand_2/b inv_2/in 0.34fF
C1462 gnd ffipg_2/ffi_1/nand_3/a 0.33fF
C1463 ffipg_3/ffi_0/inv_0/op ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C1464 ffipg_2/ffi_1/nand_7/w_0_0# ffipg_2/ffi_1/nand_7/a 0.06fF
C1465 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1466 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_6/w_0_0# 0.06fF
C1467 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_1/b 0.04fF
C1468 gnd ffipg_3/ffi_0/nand_6/a 0.37fF
C1469 ffipg_2/ffi_1/nand_1/a clk 0.13fF
C1470 sumffo_3/xor_0/inv_0/op gnd 0.32fF
C1471 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/nand_6/a 0.06fF
C1472 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C1473 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1474 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/ffo_0/nand_6/a 0.06fF
C1475 x3in clk 0.68fF
C1476 ffo_0/inv_1/w_0_6# clk 0.06fF
C1477 gnd ffipg_1/ffi_0/nand_5/w_0_0# 0.10fF
C1478 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/nand_3/b 0.06fF
C1479 sumffo_3/ffo_0/nand_1/b gnd 0.57fF
C1480 gnd sumffo_2/ffo_0/inv_0/op 0.51fF
C1481 cla_2/p0 cla_0/l 0.44fF
C1482 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/ffi_0/q 0.23fF
C1483 ffipg_2/k gnd 0.58fF
C1484 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C1485 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/nand_7/a 0.06fF
C1486 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b 0.32fF
C1487 ffipg_3/ffi_0/nand_5/w_0_0# ffipg_3/ffi_0/nand_7/a 0.04fF
C1488 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C1489 gnd ffipg_2/ffi_1/nand_4/w_0_0# 0.10fF
C1490 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# 0.04fF
C1491 sumffo_2/xor_0/inv_0/op ffi_0/q 0.06fF
C1492 gnd ffipg_3/ffi_0/nand_1/b 0.57fF
C1493 ffo_0/nand_7/a couto 0.00fF
C1494 gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C1495 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C1496 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/nand_6/a 0.06fF
C1497 ffo_0/nand_6/w_0_0# couto 0.06fF
C1498 sumffo_1/xor_0/a_10_10# gnd 0.93fF
C1499 cla_0/l cla_0/g0 0.14fF
C1500 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a 0.13fF
C1501 ffi_0/nand_1/b ffi_0/nand_7/a 0.13fF
C1502 x2in ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C1503 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/inv_1/op 0.33fF
C1504 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C1505 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C1506 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# 0.04fF
C1507 gnd sumffo_2/ffo_0/nand_7/a 0.33fF
C1508 z1o sumffo_0/ffo_0/nand_6/w_0_0# 0.06fF
C1509 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C1510 ffi_0/nand_1/a clk 0.13fF
C1511 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_3/a 0.06fF
C1512 ffipg_2/ffi_1/nand_6/w_0_0# ffipg_2/ffi_1/qbar 0.04fF
C1513 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C1514 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C1515 sumffo_2/ffo_0/nand_1/a gnd 0.33fF
C1516 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C1517 gnd nor_0/w_0_0# 0.46fF
C1518 gnd inv_7/in 0.43fF
C1519 ffo_0/qbar ffo_0/nand_6/a 0.00fF
C1520 ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1521 ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1522 ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1523 ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1524 ffipg_3/ffi_1/qbar Gnd 0.42fF
C1525 ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1526 ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1527 ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1528 ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1529 ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1530 ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1531 ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1532 ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1533 x4in Gnd 0.51fF
C1534 ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1535 ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1536 ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1537 ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1538 ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1539 ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1540 ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1541 ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1542 ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1543 ffipg_3/ffi_0/qbar Gnd 0.42fF
C1544 ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1545 ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1546 ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1547 ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1548 ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1549 ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1550 ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1551 ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1552 y4in Gnd 0.51fF
C1553 ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1554 ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1555 ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1556 ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C1557 ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1558 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1559 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1560 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1561 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1562 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1563 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1564 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1565 ffipg_3/ffi_0/q Gnd 2.68fF
C1566 ffipg_3/ffi_1/q Gnd 2.93fF
C1567 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1568 ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1569 ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1570 ffi_0/q Gnd 1.92fF
C1571 ffi_0/nand_7/a Gnd 0.30fF
C1572 ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1573 nor_0/b Gnd 1.01fF
C1574 ffi_0/nand_6/a Gnd 0.30fF
C1575 ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1576 ffi_0/inv_1/op Gnd 0.89fF
C1577 ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1578 ffi_0/nand_3/b Gnd 0.43fF
C1579 ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1580 ffi_0/nand_3/a Gnd 0.30fF
C1581 ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1582 clk Gnd 15.56fF
C1583 cinin Gnd 0.51fF
C1584 ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1585 ffi_0/inv_0/op Gnd 0.26fF
C1586 ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1587 ffi_0/nand_1/a Gnd 0.30fF
C1588 ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1589 ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1590 ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1591 ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C1592 ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1593 ffipg_2/ffi_1/qbar Gnd 0.42fF
C1594 ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C1595 ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1596 ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C1597 ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1598 ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C1599 ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1600 ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C1601 ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1602 x3in Gnd 0.51fF
C1603 ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1604 ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C1605 ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1606 ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C1607 ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1608 ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1609 ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1610 ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C1611 ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1612 ffipg_2/ffi_0/qbar Gnd 0.42fF
C1613 ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C1614 ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1615 ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C1616 ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1617 ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C1618 ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1619 ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C1620 ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1621 y3in Gnd 0.51fF
C1622 ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1623 ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C1624 ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1625 ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C1626 ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1627 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1628 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1629 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1630 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1631 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1632 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1633 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1634 ffipg_2/ffi_0/q Gnd 2.68fF
C1635 ffipg_2/ffi_1/q Gnd 2.93fF
C1636 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1637 ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1638 ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1639 ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C1640 ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1641 ffipg_1/ffi_1/qbar Gnd 0.42fF
C1642 ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C1643 ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1644 ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C1645 ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1646 ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C1647 ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1648 ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C1649 ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1650 x2in Gnd 0.51fF
C1651 ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1652 ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C1653 ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1654 ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C1655 ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1656 ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1657 ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1658 ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C1659 ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1660 ffipg_1/ffi_0/qbar Gnd 0.42fF
C1661 ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C1662 ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1663 ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C1664 ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1665 ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C1666 ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1667 ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C1668 ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1669 y2in Gnd 0.43fF
C1670 ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1671 ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C1672 ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1673 ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C1674 ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1675 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1676 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1677 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1678 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1679 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1680 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1681 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1682 ffipg_1/ffi_0/q Gnd 2.68fF
C1683 ffipg_1/ffi_1/q Gnd 2.93fF
C1684 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1685 inv_9/in Gnd 0.23fF
C1686 nor_4/w_0_0# Gnd 1.81fF
C1687 ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1688 ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1689 ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C1690 ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1691 ffipg_0/ffi_1/qbar Gnd 0.42fF
C1692 ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C1693 ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1694 ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C1695 ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1696 ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C1697 ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1698 ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C1699 ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1700 x1in Gnd 0.39fF
C1701 ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1702 ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C1703 ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1704 ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C1705 ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1706 ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1707 ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1708 ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C1709 ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1710 ffipg_0/ffi_0/qbar Gnd 0.42fF
C1711 ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C1712 ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1713 ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C1714 ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1715 ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C1716 ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1717 ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C1718 ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1719 y1in Gnd 0.51fF
C1720 ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1721 ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C1722 ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1723 ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C1724 ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1725 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1726 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1727 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1728 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1729 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1730 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1731 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1732 ffipg_0/ffi_0/q Gnd 2.68fF
C1733 ffipg_0/ffi_1/q Gnd 2.93fF
C1734 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1735 nor_4/a Gnd 0.44fF
C1736 inv_8/in Gnd 0.22fF
C1737 inv_8/w_0_6# Gnd 1.40fF
C1738 inv_7/in Gnd 0.22fF
C1739 inv_7/w_0_6# Gnd 1.40fF
C1740 inv_5/in Gnd 0.22fF
C1741 inv_5/w_0_6# Gnd 1.40fF
C1742 nor_3/b Gnd 1.17fF
C1743 cla_2/n Gnd 0.36fF
C1744 nor_4/b Gnd 0.32fF
C1745 inv_6/in Gnd 0.23fF
C1746 nor_3/w_0_0# Gnd 1.81fF
C1747 cla_1/n Gnd 0.36fF
C1748 inv_4/in Gnd 0.23fF
C1749 nor_2/w_0_0# Gnd 1.81fF
C1750 nor_2/b Gnd 1.11fF
C1751 inv_3/in Gnd 0.22fF
C1752 inv_3/w_0_6# Gnd 1.40fF
C1753 nor_1/b Gnd 0.91fF
C1754 inv_2/in Gnd 0.22fF
C1755 inv_2/w_0_6# Gnd 1.40fF
C1756 inv_1/in Gnd 0.23fF
C1757 nor_1/w_0_0# Gnd 1.81fF
C1758 inv_0/in Gnd 0.23fF
C1759 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1760 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1761 ffo_0/nand_7/a Gnd 0.30fF
C1762 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1763 ffo_0/qbar Gnd 0.42fF
C1764 ffo_0/nand_6/a Gnd 0.30fF
C1765 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1766 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1767 ffo_0/nand_3/b Gnd 0.43fF
C1768 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1769 ffo_0/nand_3/a Gnd 0.30fF
C1770 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1771 ffo_0/nand_0/b Gnd 0.63fF
C1772 ffo_0/d Gnd 0.44fF
C1773 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1774 ffo_0/inv_0/op Gnd 0.26fF
C1775 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1776 ffo_0/nand_1/a Gnd 0.30fF
C1777 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1778 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1779 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1780 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1781 ffipg_3/k Gnd 3.23fF
C1782 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1783 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1784 inv_4/op Gnd 1.37fF
C1785 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1786 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1787 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1788 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1789 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1790 sumffo_3/sbar Gnd 0.43fF
C1791 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1792 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1793 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1794 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1795 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1796 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1797 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1798 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1799 sumffo_3/ffo_0/d Gnd 0.64fF
C1800 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1801 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1802 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1803 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1804 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1805 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1806 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1807 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1808 nand_2/b Gnd 2.01fF
C1809 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1810 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1811 ffipg_1/k Gnd 3.25fF
C1812 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1813 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1814 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1815 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1816 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1817 sumffo_1/sbar Gnd 0.43fF
C1818 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1819 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1820 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1821 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1822 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1823 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1824 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1825 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1826 sumffo_1/ffo_0/d Gnd 0.64fF
C1827 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1828 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1829 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1830 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1831 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1832 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1833 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1834 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1835 ffipg_2/k Gnd 3.28fF
C1836 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1837 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1838 inv_1/op Gnd 1.37fF
C1839 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1840 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1841 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1842 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1843 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1844 sumffo_2/sbar Gnd 0.43fF
C1845 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1846 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1847 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1848 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1849 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1850 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1851 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1852 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1853 sumffo_2/ffo_0/d Gnd 0.64fF
C1854 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1855 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1856 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1857 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1858 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1859 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1860 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1861 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1862 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1863 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1864 ffipg_0/k Gnd 3.30fF
C1865 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1866 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1867 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1868 gnd Gnd 75.58fF
C1869 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1870 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1871 sumffo_0/sbar Gnd 0.43fF
C1872 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1873 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1874 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1875 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1876 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1877 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1878 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1879 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1880 sumffo_0/ffo_0/d Gnd 0.64fF
C1881 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1882 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1883 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1884 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1885 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1886 cla_2/p1 Gnd 1.09fF
C1887 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1888 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1889 cla_2/inv_0/in Gnd 0.27fF
C1890 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1891 cla_2/g1 Gnd 0.59fF
C1892 cla_2/inv_0/op Gnd 0.26fF
C1893 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1894 cla_2/p0 Gnd 1.70fF
C1895 cla_1/nor_1/w_0_0# Gnd 1.23fF
C1896 cla_1/l Gnd 0.30fF
C1897 cla_1/nor_0/w_0_0# Gnd 1.23fF
C1898 cla_1/inv_0/in Gnd 0.27fF
C1899 cla_1/inv_0/w_0_6# Gnd 0.58fF
C1900 cla_1/inv_0/op Gnd 0.26fF
C1901 cla_1/nand_0/w_0_0# Gnd 0.82fF
C1902 inv_7/op Gnd 0.26fF
C1903 cla_1/p0 Gnd 1.69fF
C1904 cla_0/nor_1/w_0_0# Gnd 1.23fF
C1905 cla_0/l Gnd 0.26fF
C1906 cla_0/nor_0/w_0_0# Gnd 1.23fF
C1907 cla_0/inv_0/in Gnd 0.27fF
C1908 cla_0/inv_0/w_0_6# Gnd 0.58fF
C1909 cla_0/inv_0/op Gnd 0.26fF
C1910 cla_0/nand_0/w_0_0# Gnd 0.82fF
C1911 cla_2/l Gnd 0.80fF
C1912 cla_0/g0 Gnd 0.70fF
C1913 inv_0/op Gnd 0.23fF
C1914 nor_0/w_0_0# Gnd 2.63fF
