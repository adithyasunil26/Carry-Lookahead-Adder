* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 gnd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 gnd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 s1 cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op s1 sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op s1 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 s1 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 s3 ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op s3 sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op s3 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 s3 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 s2 nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op s2 sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op s2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 s2 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 s4 ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op s4 sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op s4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 s4 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 gnd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 gnd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd y2in cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 cla_0/l x2in gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_0/l y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 gnd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 gnd y3in cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 cla_0/l x3in gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_0/l y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 gnd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ffipg_2/k cla_0/n 0.06fF
C1 ffipg_2/pggen_0/nand_0/w_0_0# x3in 0.06fF
C2 ffipg_3/k gnd 0.66fF
C3 cin sumffo_2/xor_0/inv_0/op 0.06fF
C4 sumffo_2/xor_0/inv_1/op inv_1/op 0.06fF
C5 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C6 cla_2/inv_0/op cla_2/nand_0/w_0_0# 0.06fF
C7 gnd inv_4/in 0.33fF
C8 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C9 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C10 nor_1/b gnd 0.35fF
C11 cla_0/g0 cla_1/p0 0.38fF
C12 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# y2in 0.23fF
C13 ffipg_3/k cla_0/l 0.10fF
C14 inv_3/w_0_6# nand_2/b 0.06fF
C15 cla_0/g0 ffipg_1/k 0.06fF
C16 y4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C17 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C18 inv_3/w_0_6# cla_1/l 0.06fF
C19 cin sumffo_0/xor_0/w_n3_4# 0.06fF
C20 sumffo_0/xor_0/inv_1/op s1 0.52fF
C21 ffipg_1/k cla_1/p0 0.05fF
C22 inv_7/w_0_6# inv_7/op 0.03fF
C23 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_0/op 0.06fF
C24 ffipg_2/pggen_0/nand_0/w_0_0# cla_2/p0 0.24fF
C25 sumffo_1/xor_0/w_n3_4# ffipg_1/k 0.06fF
C26 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C27 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C28 sumffo_2/xor_0/a_10_10# gnd 0.93fF
C29 s3 sumffo_2/xor_0/a_10_10# 0.45fF
C30 gnd inv_0/in 0.30fF
C31 x1in ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C32 gnd s2 0.14fF
C33 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C34 nor_3/b cla_2/l 0.10fF
C35 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C36 nor_3/b gnd 0.33fF
C37 cla_0/g0 cla_0/inv_0/in 0.16fF
C38 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C39 ffipg_3/k sumffo_3/xor_0/inv_0/op 0.20fF
C40 ffipg_2/k sumffo_2/xor_0/inv_0/op 0.20fF
C41 cla_2/nand_0/w_0_0# gnd 0.18fF
C42 nor_0/w_0_0# gnd 0.46fF
C43 cla_0/inv_0/in cla_1/p0 0.02fF
C44 ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.36fF
C45 cla_2/g1 cla_2/p1 0.00fF
C46 cin gnd 1.53fF
C47 cin s3 0.28fF
C48 cla_2/p1 x4in 0.22fF
C49 nor_4/w_0_0# cout 0.03fF
C50 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_1/op 0.06fF
C51 inv_1/op sumffo_2/xor_0/inv_0/op 0.27fF
C52 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C53 inv_6/in gnd 0.33fF
C54 nor_4/w_0_0# nor_4/b 0.06fF
C55 ffipg_1/pggen_0/xor_0/a_10_10# y2in 0.12fF
C56 cla_0/n inv_1/in 0.02fF
C57 sumffo_0/xor_0/inv_0/op gnd 0.36fF
C58 cla_0/inv_0/w_0_6# gnd 0.06fF
C59 nor_3/b inv_5/w_0_6# 0.17fF
C60 cin cla_0/l 0.33fF
C61 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C62 nor_2/w_0_0# inv_4/in 0.11fF
C63 gnd inv_7/in 0.43fF
C64 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C65 y3in ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C66 y4in ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C67 cin sumffo_1/xor_0/a_38_n43# 0.01fF
C68 gnd cinbar 0.16fF
C69 gnd inv_3/in 0.47fF
C70 nor_3/b nor_3/w_0_0# 0.06fF
C71 sumffo_2/xor_0/w_n3_4# gnd 0.12fF
C72 sumffo_2/xor_0/w_n3_4# s3 0.02fF
C73 gnd cla_2/n 0.60fF
C74 y3in ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C75 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C76 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/w_n3_4# 0.06fF
C77 nor_0/w_0_0# nand_2/b 0.04fF
C78 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C79 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.32fF
C80 cla_0/l inv_7/in 0.13fF
C81 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C82 cin nand_2/b 0.04fF
C83 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C84 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C85 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C86 inv_6/in nor_3/w_0_0# 0.11fF
C87 cla_1/nand_0/a_13_n26# gnd 0.01fF
C88 y1in ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C89 ffipg_0/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C90 ffipg_2/k gnd 0.64fF
C91 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C92 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C93 inv_5/in cla_0/n 0.13fF
C94 gnd y4in 1.76fF
C95 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C96 cin s4 0.16fF
C97 gnd cla_2/nor_1/w_0_0# 0.31fF
C98 gnd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C99 x3in gnd 1.24fF
C100 ffipg_0/pggen_0/xor_0/w_n3_4# y1in 0.06fF
C101 inv_1/op gnd 0.58fF
C102 cla_0/g0 nor_0/a 0.57fF
C103 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/k 0.01fF
C104 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C105 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C106 inv_8/in cin 0.13fF
C107 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C108 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C109 gnd nor_2/b 0.32fF
C110 x1in gnd 1.19fF
C111 ffipg_2/k cla_0/l 0.10fF
C112 ffipg_3/k cla_2/p1 0.05fF
C113 sumffo_0/xor_0/inv_1/op gnd 0.35fF
C114 cla_1/inv_0/in gnd 0.34fF
C115 inv_7/w_0_6# cla_2/l 0.06fF
C116 cla_1/p0 nor_0/a 0.24fF
C117 nand_2/b inv_3/in 0.13fF
C118 gnd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C119 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C120 inv_7/w_0_6# gnd 0.15fF
C121 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_0/op 0.08fF
C122 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C123 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C124 nor_3/w_0_0# cla_2/n 0.06fF
C125 ffipg_1/k nor_0/a 0.06fF
C126 gnd inv_2/in 0.47fF
C127 x1in y1in 0.73fF
C128 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C129 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C130 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C131 cin inv_8/w_0_6# 0.06fF
C132 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C133 sumffo_3/xor_0/w_n3_4# gnd 0.12fF
C134 cla_2/inv_0/in gnd 0.34fF
C135 cla_0/l cla_1/inv_0/in 0.23fF
C136 inv_0/op gnd 0.27fF
C137 cla_2/p0 cla_2/l 0.16fF
C138 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C139 inv_7/w_0_6# cla_0/l 0.06fF
C140 ffipg_2/k nand_2/b 0.06fF
C141 cla_2/p0 gnd 1.12fF
C142 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.15fF
C143 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/k 0.45fF
C144 ffipg_0/pggen_0/nand_0/w_0_0# gnd 0.10fF
C145 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C146 cla_0/nor_1/w_0_0# gnd 0.31fF
C147 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C148 gnd sumffo_3/xor_0/a_10_10# 0.93fF
C149 ffipg_0/k gnd 0.74fF
C150 cla_0/nand_0/a_13_n26# gnd 0.00fF
C151 y1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C152 gnd sumffo_1/xor_0/inv_1/op 0.35fF
C153 cla_2/inv_0/in cla_0/l 0.16fF
C154 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C155 cla_1/inv_0/op cla_0/n 0.06fF
C156 s1 sumffo_0/xor_0/w_n3_4# 0.02fF
C157 cla_2/p0 cla_0/l 0.44fF
C158 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C159 y1in ffipg_0/k 0.07fF
C160 inv_2/w_0_6# nor_1/b 0.03fF
C161 cla_0/nor_1/w_0_0# cla_0/l 0.02fF
C162 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C163 nand_2/b inv_2/in 0.34fF
C164 gnd inv_1/in 0.33fF
C165 cin sumffo_3/xor_0/a_38_n43# 0.01fF
C166 cla_0/nor_0/w_0_0# gnd 0.31fF
C167 cla_1/n inv_4/in 0.02fF
C168 ffipg_2/pggen_0/nand_0/w_0_0# gnd 0.10fF
C169 ffipg_2/pggen_0/nand_0/a_13_n26# gnd 0.01fF
C170 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# 0.16fF
C171 sumffo_2/xor_0/inv_1/op gnd 0.35fF
C172 sumffo_2/xor_0/inv_1/op s3 0.52fF
C173 cla_2/l cla_0/n 0.32fF
C174 nor_2/w_0_0# nor_2/b 0.06fF
C175 gnd cla_0/n 1.18fF
C176 cla_1/nor_0/w_0_0# gnd 0.31fF
C177 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C178 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C179 cla_2/p0 cla_1/l 0.02fF
C180 sumffo_3/xor_0/w_n3_4# s4 0.02fF
C181 ffipg_3/k inv_4/op 0.09fF
C182 s1 gnd 0.14fF
C183 inv_7/op gnd 0.27fF
C184 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C185 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C186 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C187 ffipg_2/pggen_0/nand_0/w_0_0# cla_0/l 0.04fF
C188 sumffo_3/xor_0/inv_1/w_0_6# gnd 0.06fF
C189 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C190 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C191 inv_4/op inv_4/in 0.04fF
C192 x2in y2in 0.73fF
C193 cla_2/nand_0/a_13_n26# gnd 0.01fF
C194 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C195 nor_0/w_0_0# cla_0/g0 0.06fF
C196 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C197 cla_0/l cla_0/n 0.25fF
C198 cla_2/l inv_5/in 0.05fF
C199 cla_1/nor_0/w_0_0# cla_0/l 0.01fF
C200 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C201 cin inv_2/w_0_6# 0.06fF
C202 sumffo_1/xor_0/w_n3_4# s2 0.02fF
C203 cin cla_0/g0 0.08fF
C204 s4 sumffo_3/xor_0/a_10_10# 0.45fF
C205 gnd inv_5/in 0.49fF
C206 gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C207 sumffo_3/xor_0/inv_1/op gnd 0.35fF
C208 inv_5/w_0_6# cla_0/n 0.06fF
C209 gnd sumffo_0/xor_0/inv_1/w_0_6# 0.07fF
C210 ffipg_1/pggen_0/nor_0/w_0_0# y2in 0.06fF
C211 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C212 cin ffipg_1/k 0.06fF
C213 cin sumffo_1/xor_0/w_n3_4# 0.00fF
C214 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C215 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C216 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# gnd 0.11fF
C217 nand_2/b cla_0/n 0.06fF
C218 cla_2/p1 y4in 0.03fF
C219 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C220 gnd y2in 1.82fF
C221 cla_1/l cla_0/n 0.07fF
C222 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/k 0.45fF
C223 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C224 ffipg_3/k x4in 0.46fF
C225 nor_1/b nor_1/w_0_0# 0.06fF
C226 sumffo_2/xor_0/inv_0/op gnd 0.32fF
C227 inv_5/w_0_6# inv_5/in 0.10fF
C228 s3 sumffo_2/xor_0/inv_0/op 0.06fF
C229 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C230 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C231 cla_2/inv_0/op gnd 0.27fF
C232 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# x2in 0.06fF
C233 x2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C234 cla_0/l y2in 0.13fF
C235 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C236 sumffo_0/xor_0/w_n3_4# gnd 0.12fF
C237 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C238 cla_2/inv_0/in cla_2/p1 0.02fF
C239 gnd x2in 1.24fF
C240 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C241 gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C242 ffipg_2/k cla_1/p0 0.06fF
C243 sumffo_3/xor_0/inv_1/op s4 0.52fF
C244 gnd cla_1/nor_1/w_0_0# 0.31fF
C245 cla_1/inv_0/op gnd 0.27fF
C246 cla_2/p0 cla_2/p1 0.24fF
C247 gnd ffipg_0/pggen_0/nand_0/a_13_n26# 0.01fF
C248 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C249 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C250 ffipg_1/pggen_0/xor_0/w_n3_4# y2in 0.06fF
C251 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C252 cla_1/inv_0/w_0_6# cla_1/inv_0/op 0.03fF
C253 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C254 sumffo_1/xor_0/a_10_10# s2 0.45fF
C255 inv_8/w_0_6# inv_7/op 0.06fF
C256 gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C257 gnd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C258 sumffo_1/xor_0/inv_0/op s2 0.06fF
C259 inv_2/w_0_6# inv_2/in 0.10fF
C260 cla_2/g1 cla_2/nand_0/w_0_0# 0.06fF
C261 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C262 cla_1/inv_0/op cla_0/l 0.35fF
C263 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C264 cla_1/n nor_2/b 0.39fF
C265 cla_2/l gnd 0.61fF
C266 cin sumffo_1/xor_0/a_10_10# 0.06fF
C267 cin sumffo_0/xor_0/a_10_10# 0.12fF
C268 ffipg_3/pggen_0/xor_0/inv_0/op x4in 0.27fF
C269 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C270 y3in ffipg_2/k 0.07fF
C271 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C272 s3 gnd 0.14fF
C273 sumffo_1/xor_0/inv_0/op cin 0.06fF
C274 inv_0/op cla_0/g0 0.32fF
C275 inv_6/in nor_4/b 0.04fF
C276 nor_4/a gnd 0.40fF
C277 cla_1/nand_0/w_0_0# gnd 0.10fF
C278 cla_1/inv_0/w_0_6# gnd 0.06fF
C279 x3in ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C280 y3in x3in 0.73fF
C281 y1in gnd 1.77fF
C282 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C283 nor_0/a inv_0/in 0.02fF
C284 y4in ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C285 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C286 ffipg_1/pggen_0/xor_0/w_n3_4# x2in 0.06fF
C287 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C288 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C289 cla_2/p0 cla_1/p0 0.24fF
C290 cla_2/l cla_0/l 0.37fF
C291 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C292 cla_0/l gnd 3.30fF
C293 x3in ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C294 nor_0/w_0_0# nor_0/a 0.06fF
C295 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C296 cla_2/l inv_5/w_0_6# 0.08fF
C297 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C298 inv_5/w_0_6# gnd 0.42fF
C299 cla_2/g1 cla_2/n 0.13fF
C300 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C301 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C302 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C303 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C304 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C305 sumffo_0/xor_0/inv_0/w_0_6# ffipg_0/k 0.06fF
C306 gnd nor_3/w_0_0# 0.14fF
C307 inv_9/in gnd 0.33fF
C308 ffipg_1/pggen_0/xor_0/w_n3_4# gnd 0.15fF
C309 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C310 nand_2/b gnd 1.92fF
C311 y3in cla_2/p0 0.03fF
C312 ffipg_1/pggen_0/nand_0/w_0_0# y2in 0.06fF
C313 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C314 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C315 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C316 ffipg_2/pggen_0/xor_0/a_10_10# gnd 0.93fF
C317 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C318 inv_1/op nor_1/w_0_0# 0.03fF
C319 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C320 nor_4/a inv_9/in 0.02fF
C321 cla_1/l gnd 0.40fF
C322 cla_2/g1 y4in 0.13fF
C323 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.35fF
C324 gnd sumffo_3/xor_0/inv_0/op 0.32fF
C325 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C326 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C327 x4in y4in 0.73fF
C328 nor_0/a cinbar 0.32fF
C329 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C330 gnd s4 0.14fF
C331 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C332 ffipg_1/pggen_0/xor_0/inv_0/op y2in 0.20fF
C333 y1in ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C334 cla_1/nor_0/w_0_0# cla_1/p0 0.06fF
C335 nand_2/b cla_0/l 0.06fF
C336 cla_0/l cla_1/l 0.08fF
C337 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C338 inv_8/in gnd 0.43fF
C339 nor_2/w_0_0# gnd 0.17fF
C340 sumffo_1/xor_0/inv_1/w_0_6# gnd 0.06fF
C341 inv_3/w_0_6# inv_3/in 0.10fF
C342 inv_8/in nor_4/a 0.04fF
C343 x2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C344 y3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C345 ffipg_0/pggen_0/xor_0/a_10_10# gnd 0.93fF
C346 y4in ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C347 ffipg_2/k sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C348 cla_2/inv_0/in cla_2/g1 0.04fF
C349 inv_8/w_0_6# gnd 0.15fF
C350 x4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C351 ffipg_0/pggen_0/xor_0/a_10_10# y1in 0.12fF
C352 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C353 nand_2/b cla_1/l 0.31fF
C354 cin sumffo_2/xor_0/a_38_n43# 0.01fF
C355 ffipg_1/pggen_0/xor_0/inv_0/op x2in 0.27fF
C356 nor_4/a inv_8/w_0_6# 0.03fF
C357 x1in nor_0/a 0.22fF
C358 nor_0/w_0_0# inv_0/in 0.11fF
C359 ffipg_3/pggen_0/nor_0/w_0_0# y4in 0.06fF
C360 cin sumffo_2/xor_0/a_10_10# 0.04fF
C361 cla_1/p0 y2in 0.03fF
C362 inv_1/in nor_1/w_0_0# 0.11fF
C363 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C364 cin inv_0/in 0.07fF
C365 gnd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C366 sumffo_3/xor_0/inv_0/op s4 0.06fF
C367 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C368 cin s2 0.27fF
C369 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C370 ffipg_1/k y2in 0.07fF
C371 inv_3/w_0_6# nor_2/b 0.03fF
C372 x1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C373 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C374 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C375 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C376 cin nor_0/w_0_0# 0.16fF
C377 ffipg_3/k y4in 0.07fF
C378 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C379 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.36fF
C380 nor_3/b inv_6/in 0.16fF
C381 cla_0/n nor_1/w_0_0# 0.06fF
C382 ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C383 cla_2/l cla_2/p1 0.02fF
C384 y3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C385 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C386 cla_2/p1 gnd 1.00fF
C387 y1in ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C388 cinbar inv_0/in 0.16fF
C389 ffipg_0/k nor_0/a 0.05fF
C390 nor_4/w_0_0# gnd 0.15fF
C391 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C392 cin sumffo_0/xor_0/inv_0/op 0.20fF
C393 cla_1/p0 x2in 0.22fF
C394 ffipg_1/pggen_0/xor_0/inv_1/op y2in 0.22fF
C395 nor_4/w_0_0# nor_4/a 0.07fF
C396 s1 sumffo_0/xor_0/a_10_10# 0.45fF
C397 ffipg_1/k x2in 0.46fF
C398 inv_4/in nor_2/b 0.16fF
C399 nor_0/w_0_0# cinbar 0.06fF
C400 cla_0/nand_0/w_0_0# gnd 0.10fF
C401 cla_0/l cla_2/p1 0.30fF
C402 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C403 nor_3/b cla_2/n 0.41fF
C404 inv_8/in inv_8/w_0_6# 0.10fF
C405 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C406 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C407 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C408 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C409 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C410 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C411 cin sumffo_2/xor_0/w_n3_4# 0.00fF
C412 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C413 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C414 nor_1/b inv_2/in 0.04fF
C415 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C416 inv_2/w_0_6# gnd 0.17fF
C417 ffipg_3/k cla_2/p0 0.06fF
C418 cla_0/g0 gnd 1.23fF
C419 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_1/w_0_6# 0.03fF
C420 sumffo_2/xor_0/inv_0/w_0_6# gnd 0.09fF
C421 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C422 cla_0/nand_0/w_0_0# cla_0/l 0.06fF
C423 inv_6/in cla_2/n 0.02fF
C424 cla_1/p0 gnd 1.12fF
C425 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C426 y1in cla_0/g0 0.13fF
C427 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C428 sumffo_1/xor_0/w_n3_4# gnd 0.12fF
C429 ffipg_1/k gnd 0.76fF
C430 x2in ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C431 gnd cla_1/n 0.52fF
C432 ffipg_3/pggen_0/xor_0/inv_0/op y4in 0.20fF
C433 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# x4in 0.06fF
C434 nor_4/w_0_0# inv_9/in 0.11fF
C435 inv_2/w_0_6# cla_0/l 0.06fF
C436 sumffo_0/xor_0/inv_0/w_0_6# gnd 0.11fF
C437 cla_0/g0 cla_0/l 0.14fF
C438 inv_3/w_0_6# cla_0/n 0.16fF
C439 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C440 cla_1/p0 cla_0/l 0.09fF
C441 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C442 sumffo_0/xor_0/inv_1/op cin 0.22fF
C443 cla_0/l cla_1/n 0.13fF
C444 inv_0/op inv_0/in 0.04fF
C445 cla_2/inv_0/op cla_2/g1 0.35fF
C446 ffipg_2/pggen_0/xor_0/inv_1/op gnd 0.39fF
C447 y3in gnd 1.82fF
C448 nor_1/b inv_1/in 0.16fF
C449 cla_0/inv_0/in gnd 0.34fF
C450 cin inv_2/in 0.13fF
C451 inv_2/w_0_6# nand_2/b 0.03fF
C452 inv_4/op gnd 0.58fF
C453 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C454 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C455 cla_0/g0 nand_2/b 0.13fF
C456 ffipg_3/k cla_0/n 0.06fF
C457 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.39fF
C458 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C459 sumffo_2/xor_0/w_n3_4# ffipg_2/k 0.06fF
C460 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_0/op 0.08fF
C461 cla_2/nor_0/w_0_0# gnd 0.31fF
C462 inv_0/op nor_0/w_0_0# 0.10fF
C463 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.36fF
C464 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C465 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C466 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C467 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C468 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C469 cla_1/p0 cla_1/l 0.16fF
C470 y3in cla_0/l 0.13fF
C471 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/k 0.02fF
C472 ffipg_1/k nand_2/b 0.15fF
C473 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C474 s2 sumffo_1/xor_0/inv_1/op 0.52fF
C475 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C476 nor_1/b cla_0/n 0.36fF
C477 inv_7/w_0_6# inv_7/in 0.10fF
C478 inv_3/in nor_2/b 0.04fF
C479 cla_0/inv_0/in cla_0/l 0.07fF
C480 cin sumffo_3/xor_0/a_10_10# 0.04fF
C481 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C482 cin ffipg_0/k 0.19fF
C483 cin sumffo_1/xor_0/inv_1/op 0.04fF
C484 gnd nor_1/w_0_0# 0.17fF
C485 x1in ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C486 ffipg_2/k x3in 0.46fF
C487 inv_1/op ffipg_2/k 0.09fF
C488 cout gnd 0.25fF
C489 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C490 ffipg_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C491 y3in ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C492 x1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C493 gnd nor_4/b 0.25fF
C494 cla_2/g1 gnd 0.65fF
C495 sumffo_1/xor_0/a_10_10# gnd 0.93fF
C496 sumffo_0/xor_0/a_10_10# gnd 0.93fF
C497 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C498 gnd x4in 1.24fF
C499 nor_2/w_0_0# cla_1/n 0.06fF
C500 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C501 ffipg_1/pggen_0/nand_0/a_13_n26# gnd 0.01fF
C502 nor_4/a nor_4/b 0.42fF
C503 sumffo_1/xor_0/inv_0/op gnd 0.32fF
C504 cla_2/inv_0/w_0_6# gnd 0.06fF
C505 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C506 sumffo_2/xor_0/inv_1/op cin 0.04fF
C507 ffipg_0/k cinbar 0.06fF
C508 cla_2/g1 cla_0/l 0.26fF
C509 y4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C510 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# x3in 0.06fF
C511 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C512 cla_0/inv_0/op gnd 0.27fF
C513 ffipg_2/k cla_2/p0 0.05fF
C514 cin inv_7/op 0.31fF
C515 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C516 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C517 nor_2/w_0_0# inv_4/op 0.03fF
C518 gnd nor_0/a 0.58fF
C519 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C520 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.35fF
C521 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C522 nor_3/b inv_5/in 0.04fF
C523 cla_2/p0 x3in 0.22fF
C524 gnd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C525 x3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C526 inv_9/in cout 0.04fF
C527 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/k 0.02fF
C528 sumffo_1/xor_0/inv_0/w_0_6# gnd 0.09fF
C529 s1 sumffo_0/xor_0/inv_0/op 0.06fF
C530 y1in nor_0/a 0.03fF
C531 nor_4/b nor_3/w_0_0# 0.03fF
C532 inv_9/in nor_4/b 0.16fF
C533 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C534 cla_0/inv_0/op cla_0/l 0.35fF
C535 cin sumffo_3/xor_0/inv_1/op 0.04fF
C536 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C537 cla_2/p0 cla_1/inv_0/in 0.02fF
C538 gnd ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C539 x1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C540 inv_7/op inv_7/in 0.04fF
C541 inv_3/w_0_6# gnd 0.17fF
C542 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C543 cin sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C544 cla_0/l nor_0/a 0.16fF
C545 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C546 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C547 x1in ffipg_0/k 0.46fF
C548 y1in ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C549 sumffo_0/xor_0/inv_1/op ffipg_0/k 0.06fF
C550 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C551 inv_1/op inv_1/in 0.04fF
C552 sumffo_2/xor_0/inv_1/op ffipg_2/k 0.22fF
C553 cla_0/inv_0/op nand_2/b 0.09fF
C554 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C555 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C556 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C557 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C558 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C559 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C560 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C561 y4in Gnd 2.72fF
C562 x4in Gnd 2.80fF
C563 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C564 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C565 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C566 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C567 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C568 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C569 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C570 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C571 y3in Gnd 2.72fF
C572 x3in Gnd 2.80fF
C573 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C574 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C575 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C576 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C577 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C578 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C579 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C580 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C581 y2in Gnd 2.72fF
C582 x2in Gnd 2.80fF
C583 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C584 cout Gnd 0.19fF
C585 inv_9/in Gnd 0.23fF
C586 nor_4/w_0_0# Gnd 1.81fF
C587 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C588 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C589 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C590 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C591 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C592 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C593 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C594 y1in Gnd 2.72fF
C595 x1in Gnd 2.80fF
C596 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C597 nor_4/a Gnd 0.59fF
C598 inv_8/in Gnd 0.22fF
C599 inv_8/w_0_6# Gnd 1.40fF
C600 inv_7/in Gnd 0.22fF
C601 inv_7/w_0_6# Gnd 1.40fF
C602 nor_4/b Gnd 0.32fF
C603 nor_3/b Gnd 0.77fF
C604 inv_5/in Gnd 0.22fF
C605 inv_5/w_0_6# Gnd 1.40fF
C606 cla_2/n Gnd 0.36fF
C607 inv_6/in Gnd 0.23fF
C608 nor_3/w_0_0# Gnd 1.81fF
C609 cla_1/n Gnd 0.36fF
C610 inv_4/in Gnd 0.23fF
C611 nor_2/w_0_0# Gnd 1.81fF
C612 cla_0/n Gnd 1.34fF
C613 nor_2/b Gnd 0.82fF
C614 inv_3/in Gnd 0.22fF
C615 inv_3/w_0_6# Gnd 1.40fF
C616 cinbar Gnd 1.21fF
C617 nor_0/a Gnd 2.07fF
C618 nor_1/b Gnd 1.05fF
C619 inv_2/in Gnd 0.22fF
C620 inv_2/w_0_6# Gnd 1.40fF
C621 inv_1/in Gnd 0.23fF
C622 nor_1/w_0_0# Gnd 1.81fF
C623 inv_0/in Gnd 0.23fF
C624 s4 Gnd 0.07fF
C625 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C626 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C627 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C628 ffipg_3/k Gnd 2.89fF
C629 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C630 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C631 inv_4/op Gnd 1.37fF
C632 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C633 s2 Gnd 0.07fF
C634 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C635 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C636 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C637 nand_2/b Gnd 2.33fF
C638 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C639 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C640 ffipg_1/k Gnd 2.78fF
C641 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C642 s3 Gnd 0.07fF
C643 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C644 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C645 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C646 ffipg_2/k Gnd 2.89fF
C647 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C648 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C649 inv_1/op Gnd 1.30fF
C650 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C651 s1 Gnd 0.07fF
C652 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C653 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C654 gnd Gnd 32.08fF
C655 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C656 cin Gnd 7.80fF
C657 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C658 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C659 ffipg_0/k Gnd 1.49fF
C660 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C661 cla_2/p1 Gnd 1.09fF
C662 cla_2/nor_1/w_0_0# Gnd 1.23fF
C663 cla_2/nor_0/w_0_0# Gnd 1.23fF
C664 cla_2/inv_0/in Gnd 0.27fF
C665 cla_2/inv_0/w_0_6# Gnd 0.58fF
C666 cla_2/g1 Gnd 0.59fF
C667 cla_2/inv_0/op Gnd 0.26fF
C668 cla_2/nand_0/w_0_0# Gnd 0.82fF
C669 cla_2/p0 Gnd 0.38fF
C670 cla_1/nor_1/w_0_0# Gnd 1.23fF
C671 cla_1/l Gnd 0.30fF
C672 cla_1/nor_0/w_0_0# Gnd 1.23fF
C673 cla_1/inv_0/in Gnd 0.27fF
C674 cla_1/inv_0/w_0_6# Gnd 0.58fF
C675 cla_1/inv_0/op Gnd 0.26fF
C676 cla_1/nand_0/w_0_0# Gnd 0.82fF
C677 inv_7/op Gnd 0.26fF
C678 cla_1/p0 Gnd 2.28fF
C679 cla_0/nor_1/w_0_0# Gnd 1.23fF
C680 cla_0/l Gnd 3.41fF
C681 cla_0/nor_0/w_0_0# Gnd 1.23fF
C682 cla_0/inv_0/in Gnd 0.27fF
C683 cla_0/inv_0/w_0_6# Gnd 0.58fF
C684 cla_0/inv_0/op Gnd 0.26fF
C685 cla_0/nand_0/w_0_0# Gnd 0.82fF
C686 cla_2/l Gnd 0.25fF
C687 cla_0/g0 Gnd 1.40fF
C688 inv_0/op Gnd 0.23fF
C689 nor_0/w_0_0# Gnd 2.63fF
