magic
tech scmos
timestamp 1619598025
<< error_s >>
rect 832 1038 834 1041
<< metal1 >>
rect 324 1490 391 1493
rect 396 1490 523 1493
rect 528 1490 627 1493
rect 632 1490 727 1493
rect 324 1481 561 1484
rect 558 1434 561 1481
rect 601 1460 615 1463
rect 601 1436 604 1460
rect 731 1441 733 1444
rect 324 1431 510 1434
rect 472 1328 475 1405
rect 507 1363 510 1431
rect 558 1431 599 1434
rect 558 1425 561 1431
rect 531 1406 615 1409
rect 507 1360 516 1363
rect 247 1310 249 1313
rect 513 1310 516 1360
rect 553 1348 558 1351
rect 555 1338 558 1348
rect 611 1335 617 1338
rect 652 1321 654 1324
rect 513 1307 519 1310
rect 611 1305 612 1308
rect 617 1305 642 1308
rect 472 1301 501 1304
rect 506 1301 519 1304
rect 550 1282 553 1293
rect 472 1275 494 1278
rect 499 1275 565 1278
rect 574 1276 577 1290
rect 758 1286 760 1289
rect 611 1276 620 1279
rect 248 1256 250 1259
rect 634 1251 642 1254
rect 634 1215 637 1251
rect 472 1212 637 1215
rect 472 1152 475 1212
rect 613 1181 616 1192
rect 576 1165 579 1168
rect 572 1159 579 1162
rect 637 1160 640 1163
rect 508 1149 509 1152
rect 572 1149 575 1159
rect 568 1146 575 1149
rect 247 1134 249 1137
rect 641 1134 648 1137
rect 637 1131 644 1134
rect 611 1130 637 1131
rect 472 1125 487 1128
rect 492 1125 507 1128
rect 682 1124 685 1137
rect 469 1091 472 1099
rect 501 1097 507 1100
rect 625 1092 628 1097
rect 644 1093 648 1096
rect 706 1092 714 1095
rect 469 1088 476 1091
rect 481 1088 507 1091
rect 630 1087 648 1090
rect 248 1080 250 1083
rect 706 1077 726 1080
rect 706 1076 709 1077
rect 627 1068 648 1071
rect 682 1068 685 1076
rect 830 1057 831 1060
rect 694 1038 714 1041
rect 831 1038 832 1041
rect 694 1024 697 1038
rect 472 1021 697 1024
rect 472 964 475 1021
rect 609 993 612 1004
rect 568 977 575 980
rect 570 971 575 974
rect 632 972 635 975
rect 494 961 507 964
rect 570 961 573 971
rect 568 958 573 961
rect 247 946 249 949
rect 641 946 647 949
rect 632 943 644 946
rect 609 942 633 943
rect 472 937 499 940
rect 504 937 507 940
rect 681 936 684 949
rect 469 903 472 911
rect 480 909 507 912
rect 469 900 479 903
rect 484 900 507 903
rect 625 902 628 909
rect 641 905 647 908
rect 705 904 711 907
rect 625 899 647 902
rect 248 892 250 895
rect 705 889 723 892
rect 705 888 708 889
rect 627 880 647 883
rect 681 880 684 888
rect 827 869 829 872
rect 695 850 711 853
rect 695 831 698 850
rect 472 828 698 831
rect 472 752 475 828
rect 631 793 655 796
rect 607 781 610 792
rect 631 776 634 793
rect 685 783 688 796
rect 715 783 718 797
rect 752 784 755 797
rect 709 780 718 783
rect 648 769 651 772
rect 568 765 573 768
rect 645 765 651 766
rect 567 759 573 762
rect 648 763 651 765
rect 709 764 718 767
rect 567 749 570 759
rect 565 746 570 749
rect 247 734 249 737
rect 709 735 718 738
rect 752 735 755 736
rect 685 734 688 735
rect 631 731 638 734
rect 607 730 631 731
rect 472 725 504 728
rect 672 721 675 734
rect 696 718 705 721
rect 739 708 742 721
rect 469 691 472 699
rect 484 697 504 700
rect 469 688 504 691
rect 622 687 625 697
rect 782 695 787 698
rect 634 690 638 693
rect 696 689 702 692
rect 622 684 638 687
rect 248 680 250 683
rect 699 680 702 689
rect 699 677 705 680
rect 782 679 785 695
rect 763 676 785 679
rect 607 645 610 668
rect 621 665 638 668
rect 672 665 675 673
rect 693 655 696 673
rect 693 652 705 655
rect 739 652 742 660
rect 268 642 297 645
rect 302 642 799 645
<< m2contact >>
rect 472 1405 477 1410
rect 557 1420 562 1425
rect 526 1406 531 1411
rect 647 1320 652 1325
rect 612 1304 617 1309
rect 501 1299 506 1304
rect 575 1298 580 1303
rect 494 1274 499 1279
rect 565 1275 570 1280
rect 620 1276 625 1281
rect 571 1165 576 1170
rect 640 1160 645 1165
rect 503 1149 508 1154
rect 487 1123 492 1128
rect 496 1097 501 1102
rect 639 1093 644 1098
rect 476 1087 481 1092
rect 625 1087 630 1092
rect 563 977 568 982
rect 489 961 494 966
rect 635 970 640 975
rect 499 935 504 940
rect 475 909 480 914
rect 479 898 484 903
rect 636 905 641 910
rect 607 776 612 781
rect 563 765 568 770
rect 629 760 634 765
rect 499 749 504 754
rect 479 697 484 702
rect 629 690 634 695
rect 605 668 610 673
<< metal2 >>
rect 477 1407 526 1410
rect 477 914 480 1087
rect 489 966 492 1123
rect 496 1102 499 1274
rect 503 1154 506 1299
rect 519 1195 522 1351
rect 558 1168 561 1420
rect 648 1325 651 1364
rect 622 1321 647 1324
rect 575 1280 578 1298
rect 570 1277 578 1280
rect 612 1201 615 1304
rect 622 1281 625 1321
rect 601 1198 615 1201
rect 558 1165 571 1168
rect 519 1007 522 1054
rect 601 1031 604 1198
rect 640 1098 643 1160
rect 563 1028 604 1031
rect 563 982 566 1028
rect 627 1015 630 1087
rect 579 1012 630 1015
rect 481 702 484 898
rect 501 754 504 935
rect 520 862 523 866
rect 517 859 523 862
rect 517 795 520 859
rect 579 806 582 1012
rect 636 910 639 970
rect 563 803 582 806
rect 563 770 566 803
rect 609 781 612 880
rect 607 673 610 776
rect 629 695 632 760
<< m123contact >>
rect 391 1490 396 1495
rect 523 1490 528 1495
rect 627 1490 632 1495
rect 599 1431 604 1436
rect 522 1348 527 1353
rect 647 1364 652 1369
rect 617 1334 622 1339
rect 599 1274 604 1279
rect 546 1146 551 1151
rect 613 1176 618 1181
rect 701 1121 706 1126
rect 611 1066 616 1071
rect 609 988 614 993
rect 700 933 705 938
rect 609 880 614 885
rect 559 746 564 751
rect 643 769 648 774
rect 713 770 718 775
rect 773 765 778 770
rect 643 760 648 765
rect 700 669 705 674
rect 297 640 302 645
<< metal3 >>
rect 392 1342 395 1490
rect 524 1353 527 1490
rect 628 1432 631 1490
rect 601 1357 604 1431
rect 647 1369 650 1423
rect 734 1357 737 1359
rect 601 1354 737 1357
rect 622 1335 634 1338
rect 298 1246 307 1249
rect 304 1073 307 1246
rect 298 1070 307 1073
rect 283 883 295 886
rect 304 885 307 1070
rect 283 720 286 883
rect 298 882 307 885
rect 441 732 444 1313
rect 631 1277 634 1335
rect 631 1274 654 1277
rect 600 1208 603 1274
rect 600 1205 616 1208
rect 613 1181 616 1205
rect 734 1185 737 1354
rect 734 1182 809 1185
rect 548 1103 551 1146
rect 548 1100 600 1103
rect 597 812 600 1100
rect 613 1071 616 1176
rect 706 1123 726 1126
rect 611 993 614 1066
rect 610 885 613 988
rect 705 934 723 937
rect 806 823 809 1182
rect 713 820 809 823
rect 597 809 646 812
rect 643 774 646 809
rect 713 775 716 820
rect 643 749 646 760
rect 564 746 646 749
rect 778 729 781 768
rect 702 726 781 729
rect 702 674 705 726
rect 297 645 300 670
use sumffo  sumffo_0
timestamp 1619451829
transform 1 0 618 0 -1 1503
box -3 24 113 129
use ffipg  ffipg_0
timestamp 1619450786
transform 1 0 2 0 1 1158
box 247 76 470 193
use nor  nor_0
timestamp 1618580541
transform 1 0 519 0 1 1312
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 553 0 1 1305
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 577 0 1 1311
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1619451829
transform 1 0 645 0 -1 1348
box -3 24 113 129
use ffipg  ffipg_1
timestamp 1619450786
transform 1 0 2 0 1 982
box 247 76 470 193
use nand  nand_1
timestamp 1618580231
transform 1 0 579 0 -1 1157
box 0 -35 34 27
use inv  inv_2
timestamp 1618579805
transform 1 0 613 0 -1 1164
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 1100
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 648 0 1 1098
box 0 -30 34 39
use inv  inv_1
timestamp 1618579805
transform 1 0 682 0 1 1091
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1619451829
transform 1 0 717 0 1 998
box -3 24 113 129
use ffipg  ffipg_2
timestamp 1619450786
transform 1 0 2 0 1 794
box 247 76 470 193
use nand  nand_2
timestamp 1618580231
transform 1 0 575 0 -1 969
box 0 -35 34 27
use inv  inv_3
timestamp 1618579805
transform 1 0 609 0 -1 976
box 0 -15 24 33
use cla  cla_1
timestamp 1618627066
transform 1 0 516 0 1 912
box -9 -46 112 95
use nor  nor_2
timestamp 1618580541
transform 1 0 647 0 1 910
box 0 -30 34 39
use inv  inv_4
timestamp 1618579805
transform 1 0 681 0 1 903
box 0 -15 24 33
use sumffo  sumffo_3
timestamp 1619451829
transform 1 0 714 0 1 810
box -3 24 113 129
use ffipg  ffipg_3
timestamp 1619450786
transform 1 0 2 0 1 582
box 247 76 470 193
use nand  nand_3
timestamp 1618580231
transform 1 0 573 0 -1 757
box 0 -35 34 27
use inv  inv_5
timestamp 1618579805
transform 1 0 607 0 -1 764
box 0 -15 24 33
use nand  nand_4
timestamp 1618580231
transform 1 0 651 0 -1 761
box 0 -35 34 27
use inv  inv_7
timestamp 1618579805
transform 1 0 685 0 -1 768
box 0 -15 24 33
use nand  nand_5
timestamp 1618580231
transform 1 0 718 0 -1 762
box 0 -35 34 27
use inv  inv_8
timestamp 1618579805
transform 1 0 752 0 -1 769
box 0 -15 24 33
use cla  cla_2
timestamp 1618627066
transform 1 0 513 0 1 700
box -9 -46 112 95
use nor  nor_3
timestamp 1618580541
transform 1 0 638 0 1 695
box 0 -30 34 39
use inv  inv_6
timestamp 1618579805
transform 1 0 672 0 1 688
box 0 -15 24 33
use nor  nor_4
timestamp 1618580541
transform 1 0 705 0 1 682
box 0 -30 34 39
use inv  inv_9
timestamp 1618579805
transform 1 0 739 0 1 675
box 0 -15 24 33
<< labels >>
rlabel metal1 324 1431 324 1434 1 cinbar
rlabel metal1 733 1441 733 1444 1 s1
rlabel metal1 324 1481 324 1484 1 cin
rlabel metal1 506 1491 506 1491 5 vdd!
rlabel metal1 832 1038 832 1041 7 s3
rlabel metal1 247 1310 247 1313 3 x1in
rlabel metal1 248 1256 248 1259 3 y1in
rlabel metal1 760 1286 760 1289 1 s2
rlabel metal1 247 1134 247 1137 3 x2in
rlabel metal1 248 1080 248 1083 3 y2in
rlabel metal1 247 946 247 949 3 x3in
rlabel metal1 248 892 248 895 3 y3in
rlabel metal1 829 869 829 872 7 s4
rlabel metal1 247 734 247 737 3 x4in
rlabel metal1 248 680 248 683 3 y4in
rlabel metal1 787 695 787 698 1 cout
rlabel metal1 311 643 311 643 1 gnd!
<< end >>
