* SPICE3 file created from nand.ext - technology: scmos
.include ../TSMC_180nm.txt
* D G S B
.param SUPPLY=1.8V
.param LAMBDA=0.09u
.param length={2*LAMBDA}
.param w={6*LAMBDA}
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

va a gnd pulse 1.8 0 0ns 10ps 10ps 10ns 20ns
vb b gnd pulse 1.8 0 0ns 10ps 10ps 20ns 40ns

M1000 a_13_n26# a gnd Gnd CMOSN w=12 l=2
+  ad=96 pd=40 as=60 ps=34
M1001 vdd b out w_0_0# CMOSP w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1002 out a vdd w_0_0# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out b a_13_n26# Gnd CMOSN w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 b a 0.21fF
C1 w_0_0# a 0.06fF
C2 out b 0.13fF
C3 w_0_0# out 0.04fF
C4 w_0_0# vdd 0.07fF
C5 w_0_0# b 0.06fF
C6 gnd Gnd 0.11fF
C7 out Gnd 0.07fF
C8 vdd Gnd 0.06fF
C9 b Gnd 0.20fF
C10 a Gnd 0.17fF
C11 w_0_0# Gnd 0.82fF

.tran 100p 40n

.control
set hcopypscolor = 1 
set color0=white 
set color1=black 

run
set curplottitle="Adithya-2019102005-nand"

hardcopy nand.eps v(out) 
hardcopy a.eps v(a) 
hardcopy b.eps v(b)
.endc