* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 a_33_8# a_29_2# op w_n3_2# pfet w=24 l=2
+  ad=144 pd=60 as=312 ps=74
M1005 gnd a_38_n5# a_33_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=72 ps=36
M1006 vdd a_38_n5# a_33_8# w_n3_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_10_8# a_5_n13# vdd w_n3_2# pfet w=24 l=2
+  ad=144 pd=60 as=0 ps=0
M1008 a_10_n33# a_5_n13# gnd Gnd nfet w=12 l=2
+  ad=72 pd=36 as=0 ps=0
M1009 op a_14_2# a_10_8# w_n3_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 op a_14_n20# a_10_n33# Gnd nfet w=12 l=2
+  ad=156 pd=50 as=0 ps=0
M1011 a_33_n33# a_30_n20# op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
C0 inv_1/op a_14_2# 0.03fF
C1 vdd inv_1/op 0.15fF
C2 a gnd 0.54fF
C3 m2_n10_n50# vdd 0.02fF
C4 m3_n10_n50# a 0.03fF
C5 a_30_n20# a_38_n5# 0.04fF
C6 op gnd 0.04fF
C7 m2_n18_10# inv_0/op 0.02fF
C8 w_n3_2# a_5_n13# 0.06fF
C9 inv_1/w_0_6# inv_1/in 0.06fF
C10 m3_n18_10# a_5_n13# 0.00fF
C11 inv_0/w_0_6# a 0.06fF
C12 m3_n10_n50# vdd 0.07fF
C13 m3_n18_10# a 0.04fF
C14 op w_n3_2# 0.02fF
C15 m3_n18_10# op 0.01fF
C16 w_n3_2# a_14_2# 0.08fF
C17 b inv_1/in 0.05fF
C18 a a_5_n13# 0.04fF
C19 vdd w_n3_2# 0.14fF
C20 inv_0/op gnd 0.10fF
C21 inv_0/w_0_6# vdd 0.06fF
C22 a_30_n20# inv_1/op 0.03fF
C23 m1_38_n5# a_38_n5# 0.04fF
C24 w_n3_2# a_29_2# 0.08fF
C25 a_5_n13# a_14_2# 0.04fF
C26 inv_1/w_0_6# inv_1/op 0.03fF
C27 inv_0/w_0_6# inv_0/op 0.03fF
C28 a vdd 0.02fF
C29 m3_n18_10# inv_0/op 0.02fF
C30 op vdd 0.03fF
C31 b inv_1/op 0.40fF
C32 inv_1/in inv_1/op 0.04fF
C33 a inv_0/op 0.04fF
C34 a_14_n20# a_5_n13# 0.04fF
C35 b m2_38_n5# 0.01fF
C36 m2_38_n5# a_38_n5# 0.00fF
C37 b gnd 0.16fF
C38 inv_1/in gnd 0.05fF
C39 m3_n10_n50# b 0.03fF
C40 vdd inv_0/op 0.15fF
C41 m1_38_n5# m2_38_n5# 0.01fF
C42 b w_n3_2# 0.08fF
C43 m3_n10_n50# m2_n10_36# 0.01fF
C44 a_38_n5# w_n3_2# 0.06fF
C45 m3_n18_10# b 0.04fF
C46 m3_n18_10# a_38_n5# 0.01fF
C47 b a_5_n13# 0.00fF
C48 inv_1/op gnd 0.29fF
C49 b a 0.06fF
C50 m3_n18_10# m1_38_n5# 0.00fF
C51 a inv_1/in 0.01fF
C52 vdd inv_1/w_0_6# 0.06fF
C53 m3_n10_n50# inv_1/op 0.04fF
C54 b op 0.22fF
C55 m2_n10_n50# m3_n10_n50# 0.01fF
C56 op a_38_n5# 0.06fF
C57 m3_n18_10# m2_n18_10# 0.02fF
C58 inv_1/op w_n3_2# 0.08fF
C59 vdd inv_1/in 0.02fF
C60 m3_n18_10# inv_1/op 0.25fF
C61 m3_n10_n50# gnd 0.01fF
C62 m1_38_n5# op 0.07fF
C63 m2_n10_36# vdd 0.04fF
C64 b a_29_2# 0.03fF
C65 m3_n18_10# m2_38_n5# 0.02fF
C66 a_38_n5# a_29_2# 0.04fF
C67 inv_1/op a_5_n13# 0.00fF
C68 a inv_1/op 0.16fF
C69 m3_n18_10# gnd 0.01fF
C70 b a_14_n20# 0.03fF
C71 m3_n10_n50# m3_n18_10# 0.07fF
C72 op inv_1/op 0.20fF
C73 m3_n18_10# Gnd 0.07fF **FLOATING
C74 m3_n10_n50# Gnd 0.37fF **FLOATING
C75 m2_n10_n50# Gnd 0.09fF **FLOATING
C76 m2_38_n5# Gnd 0.08fF **FLOATING
C77 m2_n18_10# Gnd 0.09fF **FLOATING
C78 m2_n10_36# Gnd 0.07fF **FLOATING
C79 m1_38_n5# Gnd 0.02fF **FLOATING
C80 b Gnd 0.88fF **FLOATING
C81 a_30_n20# Gnd 0.09fF
C82 a_14_n20# Gnd 0.09fF
C83 op Gnd 0.11fF
C84 a_38_n5# Gnd 0.19fF
C85 a_29_2# Gnd 0.01fF
C86 a_14_2# Gnd 0.01fF
C87 a_5_n13# Gnd 0.19fF
C88 w_n3_2# Gnd 1.01fF
C89 gnd Gnd 0.54fF
C90 inv_1/op Gnd 0.30fF
C91 inv_1/in Gnd 0.14fF
C92 inv_1/w_0_6# Gnd 0.58fF
C93 inv_0/op Gnd 0.08fF
C94 vdd Gnd 0.28fF
C95 a Gnd 0.98fF
C96 inv_0/w_0_6# Gnd 0.58fF
