magic
tech scmos
timestamp 1618580541
<< nwell >>
rect 0 0 34 36
<< ntransistor >>
rect 11 -21 13 -15
rect 21 -21 23 -15
<< ptransistor >>
rect 11 6 13 30
rect 21 6 23 30
<< ndiffusion >>
rect 10 -21 11 -15
rect 13 -21 15 -15
rect 19 -21 21 -15
rect 23 -21 24 -15
<< pdiffusion >>
rect 10 6 11 30
rect 13 6 21 30
rect 23 6 24 30
<< ndcontact >>
rect 6 -21 10 -15
rect 15 -21 19 -15
rect 24 -21 28 -15
<< pdcontact >>
rect 6 6 10 30
rect 24 6 28 30
<< polysilicon >>
rect 11 30 13 33
rect 21 30 23 33
rect 11 -15 13 6
rect 21 -15 23 6
rect 11 -24 13 -21
rect 21 -24 23 -21
<< polycontact >>
rect 7 -12 11 -8
rect 17 -5 21 -1
<< metal1 >>
rect 0 36 34 39
rect 6 30 9 36
rect 0 -5 17 -2
rect 25 -3 28 6
rect 25 -6 34 -3
rect 0 -11 7 -8
rect 25 -9 28 -6
rect 16 -12 28 -9
rect 16 -15 19 -12
rect 6 -27 9 -21
rect 25 -27 28 -21
rect 0 -30 34 -27
<< labels >>
rlabel metal1 18 37 18 37 5 vdd!
rlabel metal1 34 -6 34 -3 7 out
rlabel metal1 21 -28 21 -28 1 gnd!
rlabel metal1 0 -5 0 -2 3 b
rlabel metal1 0 -11 0 -8 3 a
<< end >>
