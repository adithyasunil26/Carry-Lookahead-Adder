magic
tech scmos
timestamp 1618371503
<< nwell >>
rect 0 0 34 36
<< ntransistor >>
rect 11 -19 13 -13
rect 21 -19 23 -13
<< ptransistor >>
rect 11 6 13 30
rect 21 6 23 30
<< ndiffusion >>
rect 6 -15 11 -13
rect 10 -19 11 -15
rect 13 -17 15 -13
rect 19 -17 21 -13
rect 13 -19 21 -17
rect 23 -15 28 -13
rect 23 -19 24 -15
<< pdiffusion >>
rect 10 26 11 30
rect 6 6 11 26
rect 13 6 21 30
rect 23 10 28 30
rect 23 6 24 10
<< ndcontact >>
rect 6 -19 10 -15
rect 15 -17 19 -13
rect 24 -19 28 -15
<< pdcontact >>
rect 6 26 10 30
rect 24 6 28 10
<< polysilicon >>
rect 11 30 13 33
rect 21 30 23 33
rect 11 -13 13 6
rect 21 -13 23 6
rect 11 -22 13 -19
rect 21 -22 23 -19
<< polycontact >>
rect 7 -10 11 -6
rect 17 -4 21 0
<< metal1 >>
rect 0 36 34 39
rect 6 30 9 36
rect 25 0 28 6
rect 0 -3 17 0
rect 25 -3 34 0
rect 0 -9 7 -6
rect 25 -7 28 -3
rect 16 -10 28 -7
rect 16 -13 19 -10
rect 6 -25 9 -19
rect 25 -25 28 -19
rect 0 -28 34 -25
<< labels >>
rlabel metal1 21 -26 21 -26 1 gnd!
rlabel metal1 18 37 18 37 5 vdd!
rlabel metal1 0 -3 0 0 3 b
rlabel metal1 0 -9 0 -6 3 a
rlabel metal1 34 -3 34 0 7 out
<< end >>
