magic
tech scmos
timestamp 1618500630
<< error_s >>
rect 25 -8 26 -2
<< nwell >>
rect -6 2 46 38
<< ntransistor >>
rect 5 -33 7 -21
rect 12 -33 14 -21
rect 26 -33 28 -21
rect 33 -33 35 -21
<< ptransistor >>
rect 5 8 7 32
rect 12 8 14 32
rect 26 8 28 32
rect 33 8 35 32
<< ndiffusion >>
rect 0 -29 5 -21
rect 4 -33 5 -29
rect 7 -33 12 -21
rect 14 -25 18 -21
rect 22 -25 26 -21
rect 14 -33 26 -25
rect 28 -33 33 -21
rect 35 -29 40 -21
rect 35 -33 36 -29
<< pdiffusion >>
rect 4 28 5 32
rect 0 8 5 28
rect 7 8 12 32
rect 14 12 26 32
rect 14 8 18 12
rect 22 8 26 12
rect 28 8 33 32
rect 35 28 36 32
rect 35 8 40 28
<< ndcontact >>
rect 0 -33 4 -29
rect 18 -25 22 -21
rect 36 -33 40 -29
<< pdcontact >>
rect 0 28 4 32
rect 18 8 22 12
rect 36 28 40 32
<< polysilicon >>
rect 5 32 7 35
rect 12 32 14 35
rect 26 32 28 35
rect 33 32 35 35
rect 5 -21 7 8
rect 12 7 14 8
rect 26 7 28 8
rect 11 3 15 7
rect 25 -20 30 -15
rect 12 -21 14 -20
rect 26 -21 28 -20
rect 33 -21 35 8
rect 5 -36 7 -33
rect 12 -36 14 -33
rect 26 -36 28 -33
rect 33 -36 35 -33
<< polycontact >>
rect 1 -12 5 -8
rect 25 3 29 7
rect 29 -5 33 -1
rect 11 -20 15 -16
<< metal1 >>
rect -15 38 46 41
rect 0 32 3 38
rect 37 32 40 38
rect -51 10 -50 13
rect -15 10 -10 15
rect 19 -8 22 8
rect 19 -11 46 -8
rect -51 -21 -50 -18
rect -19 -19 -12 -18
rect -15 -23 -12 -19
rect 19 -21 22 -11
rect 0 -37 3 -33
rect 37 -37 40 -33
rect -6 -40 46 -37
<< m2contact >>
rect -50 9 -45 14
rect -50 -22 -45 -17
<< metal2 >>
rect -15 10 -10 15
rect -49 1 -46 9
rect 25 3 29 7
rect -49 -2 -10 1
rect -13 -8 -10 -2
rect 15 -8 22 -6
rect 25 -8 28 3
rect -13 -11 5 -8
rect -48 -14 -17 -11
rect 1 -12 5 -11
rect 12 -11 28 -8
rect -48 -17 -45 -14
rect -20 -15 -17 -14
rect -20 -16 -9 -15
rect 12 -16 15 -11
rect -20 -17 -3 -16
rect 11 -17 15 -16
rect -20 -18 15 -17
rect -12 -19 15 -18
rect -6 -20 15 -19
<< m123contact >>
rect 10 2 15 7
rect 25 -20 30 -15
rect -15 -28 -10 -23
<< metal3 >>
rect 12 -5 15 2
rect -6 -6 15 -5
rect -6 -8 28 -6
rect -6 -24 -3 -8
rect 12 -9 28 -8
rect 25 -15 28 -9
rect -10 -27 -3 -24
<< metal4 >>
rect -13 -2 -10 10
rect 29 -2 33 -1
rect -13 -5 33 -2
<< m345contact >>
rect -15 10 -10 15
use inv  inv_0
timestamp 1618367270
transform 1 0 -42 0 1 8
box -3 -13 27 33
use inv  inv_1
timestamp 1618367270
transform 1 0 -42 0 -1 -15
box -3 -13 27 33
<< labels >>
rlabel metal1 -51 -21 -51 -18 3 b
rlabel metal1 -51 10 -51 13 3 a
rlabel metal1 46 -11 46 -8 7 op
rlabel metal1 20 40 20 40 5 vdd!
rlabel metal1 21 -39 21 -39 1 gnd!
<< end >>
