* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 vdd a_35_n5# a_30_8# w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=144 ps=60
M1005 a_7_8# a vdd w_n6_2# pfet w=24 l=2
+  ad=144 pd=60 as=0 ps=0
M1006 a_30_n33# a_27_n20# op Gnd nfet w=12 l=2
+  ad=72 pd=36 as=156 ps=50
M1007 op a_11_2# a_7_8# w_n6_2# pfet w=24 l=2
+  ad=312 pd=74 as=0 ps=0
M1008 gnd a_35_n5# a_30_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_7_n33# a gnd Gnd nfet w=12 l=2
+  ad=72 pd=36 as=0 ps=0
M1010 op b a_7_n33# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_30_8# b op w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 op m1_35_n5# 0.07fF
C1 inv_0/op a 0.08fF
C2 a_35_n5# a_27_n20# 0.04fF
C3 inv_1/op op 0.20fF
C4 vdd b 0.03fF
C5 inv_0/op inv_0/w_0_6# 0.04fF
C6 b gnd 0.13fF
C7 vdd a 0.03fF
C8 a gnd 0.42fF
C9 m2_n15_10# inv_0/op 0.02fF
C10 inv_1/op a_27_n20# 0.03fF
C11 a b 0.11fF
C12 vdd inv_0/w_0_6# 0.06fF
C13 op w_n6_2# 0.02fF
C14 m3_n15_10# op 0.01fF
C15 a_35_n5# b 0.04fF
C16 a inv_0/w_0_6# 0.08fF
C17 inv_1/op vdd 0.15fF
C18 inv_1/op gnd 0.12fF
C19 m3_n15_10# inv_0/op 0.02fF
C20 a_35_n5# m1_35_n5# 0.04fF
C21 a a_11_2# 0.04fF
C22 inv_1/op b 0.44fF
C23 inv_1/op a 0.15fF
C24 vdd w_n6_2# 0.09fF
C25 m2_35_n5# b 0.01fF
C26 b w_n6_2# 0.16fF
C27 a w_n6_2# 0.06fF
C28 m3_n15_10# b 0.04fF
C29 m3_n15_10# a 0.04fF
C30 a_35_n5# m2_35_n5# 0.00fF
C31 a_35_n5# w_n6_2# 0.06fF
C32 inv_1/w_0_6# vdd 0.06fF
C33 inv_1/op a_11_2# 0.03fF
C34 m2_35_n5# m1_35_n5# 0.01fF
C35 a_35_n5# m3_n15_10# 0.01fF
C36 m3_n15_10# m1_35_n5# 0.00fF
C37 m3_n15_10# m2_n15_10# 0.02fF
C38 inv_1/w_0_6# b 0.08fF
C39 a_11_2# w_n6_2# 0.08fF
C40 inv_1/op w_n6_2# 0.08fF
C41 inv_1/op m3_n15_10# 0.25fF
C42 op b 0.22fF
C43 m3_n15_10# m2_35_n5# 0.02fF
C44 inv_0/op vdd 0.15fF
C45 inv_0/op gnd 0.12fF
C46 a_35_n5# op 0.06fF
C47 inv_1/op inv_1/w_0_6# 0.04fF
C48 m3_n15_10# Gnd 0.11fF **FLOATING
C49 m2_35_n5# Gnd 0.08fF **FLOATING
C50 m2_n15_10# Gnd 0.09fF **FLOATING
C51 m1_35_n5# Gnd 0.02fF **FLOATING
C52 a_27_n20# Gnd 0.09fF
C53 op Gnd 0.14fF
C54 a_35_n5# Gnd 0.19fF
C55 a_11_2# Gnd 0.01fF
C56 w_n6_2# Gnd 1.99fF
C57 gnd Gnd 0.39fF
C58 inv_1/op Gnd 0.38fF
C59 b Gnd 1.41fF
C60 inv_1/w_0_6# Gnd 0.58fF
C61 inv_0/op Gnd 0.08fF
C62 vdd Gnd 0.23fF
C63 a Gnd 1.10fF
C64 inv_0/w_0_6# Gnd 0.58fF
