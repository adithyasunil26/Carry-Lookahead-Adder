* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=180 ps=112
M1001 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1002 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 a_7_8# a_1_n12# vdd w_n6_2# pfet w=24 l=2
+  ad=120 pd=58 as=0 ps=0
M1005 a_28_8# a_25_3# op w_n6_2# pfet w=24 l=2
+  ad=120 pd=58 as=288 ps=72
M1006 op a_11_3# a_7_8# w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_n32# a_1_n12# gnd Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 op a_11_n19# a_7_n32# Gnd nfet w=12 l=2
+  ad=144 pd=48 as=0 ps=0
M1009 a_28_n32# a_25_n19# op Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1010 gnd a_29_n5# a_28_n32# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 vdd a_29_n5# a_28_8# w_n6_2# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 inv_1/op a_25_n19# 0.01fF
C1 b a 0.07fF
C2 inv_1/w_0_6# vdd 0.06fF
C3 a_25_n19# a_29_n5# 0.04fF
C4 inv_1/op vdd 0.15fF
C5 gnd a 0.42fF
C6 m3_n15_10# op 0.00fF
C7 m3_n15_10# b 0.10fF
C8 w_n6_2# a_25_3# 0.09fF
C9 inv_1/op a 0.12fF
C10 op a_25_3# 0.05fF
C11 b a_25_3# 0.02fF
C12 m2_n15_10# inv_0/op 0.02fF
C13 inv_0/op vdd 0.15fF
C14 a_1_n12# w_n6_2# 0.06fF
C15 m3_n15_10# inv_1/op 0.24fF
C16 m3_n15_10# a_29_n5# 0.00fF
C17 a_1_n12# b 0.00fF
C18 inv_0/op a 0.08fF
C19 a_1_n12# a_11_3# 0.04fF
C20 a_29_n5# a_25_3# 0.04fF
C21 m3_n15_10# inv_0/op 0.02fF
C22 vdd a 0.03fF
C23 inv_0/op inv_0/w_0_6# 0.04fF
C24 a_1_n12# inv_1/op 0.02fF
C25 w_n6_2# op 0.02fF
C26 w_n6_2# b 0.07fF
C27 m2_n15_10# m3_n15_10# 0.02fF
C28 vdd inv_0/w_0_6# 0.06fF
C29 b op 0.12fF
C30 w_n6_2# a_11_3# 0.09fF
C31 gnd b 0.13fF
C32 op a_11_3# 0.04fF
C33 m3_n15_10# a 0.04fF
C34 a inv_0/w_0_6# 0.08fF
C35 b inv_1/w_0_6# 0.08fF
C36 w_n6_2# inv_1/op 0.00fF
C37 w_n6_2# a_29_n5# 0.06fF
C38 inv_1/op op 0.08fF
C39 inv_1/op b 0.34fF
C40 op a_29_n5# 0.14fF
C41 a_1_n12# a_11_n19# 0.04fF
C42 gnd inv_1/op 0.12fF
C43 inv_1/op a_11_3# 0.01fF
C44 a_1_n12# a 0.02fF
C45 inv_1/op inv_1/w_0_6# 0.04fF
C46 a_25_n19# op 0.10fF
C47 m3_n15_10# a_1_n12# 0.00fF
C48 w_n6_2# vdd 0.09fF
C49 gnd inv_0/op 0.12fF
C50 b vdd 0.03fF
C51 a_11_n19# op 0.04fF
C52 a_11_n19# b 0.04fF
C53 m3_n15_10# Gnd 0.07fF **FLOATING
C54 m2_n15_10# Gnd 0.09fF **FLOATING
C55 a_25_n19# Gnd 0.09fF
C56 a_11_n19# Gnd 0.09fF
C57 op Gnd 0.13fF
C58 a_29_n5# Gnd 0.20fF
C59 a_1_n12# Gnd 0.20fF
C60 w_n6_2# Gnd 1.88fF
C61 gnd Gnd 0.38fF
C62 inv_1/op Gnd 0.22fF
C63 b Gnd 1.27fF
C64 inv_1/w_0_6# Gnd 0.58fF
C65 inv_0/op Gnd 0.08fF
C66 vdd Gnd 0.23fF
C67 a Gnd 0.88fF
C68 inv_0/w_0_6# Gnd 0.58fF
