magic
tech scmos
timestamp 1618623899
<< metal1 >>
rect -4 237 0 240
rect 216 207 231 210
rect -3 156 0 187
rect 221 173 224 181
rect -4 153 0 156
rect -3 83 0 153
rect 221 89 224 98
rect 228 79 231 207
rect 469 170 470 173
rect 247 152 249 155
rect 469 143 470 146
rect 469 117 470 120
rect 247 98 249 101
rect 228 76 243 79
rect 228 63 231 76
rect 215 60 231 63
rect -4 30 0 33
<< m2contact >>
rect 219 168 224 173
rect 219 98 224 103
rect 242 151 247 156
rect 242 98 247 103
<< metal2 >>
rect 221 155 224 168
rect 221 152 242 155
rect 224 98 242 101
<< m123contact >>
rect 173 266 178 271
rect 261 182 266 187
rect 173 146 178 151
rect 173 119 178 124
rect 293 88 298 93
rect 243 76 248 81
rect 173 1 178 6
<< metal3 >>
rect 170 148 173 269
rect 237 182 261 185
rect 174 136 177 146
rect 237 136 240 182
rect 174 133 240 136
rect 174 124 177 133
rect 170 1 173 122
rect 293 81 296 88
rect 248 78 296 81
use ffi  ffi_1
timestamp 1618618094
transform 1 0 14 0 1 179
box -14 -42 207 91
use ffi  ffi_0
timestamp 1618618094
transform 1 0 14 0 -1 91
box -14 -42 207 91
use pggen  pggen_0
timestamp 1618621484
transform 1 0 250 0 1 82
box -1 -6 219 111
<< labels >>
rlabel metal1 -4 30 -4 33 3 y
rlabel metal1 -4 237 -4 240 3 x
rlabel metal1 -4 153 -4 156 3 clk
rlabel metal1 470 170 470 173 7 k
rlabel metal1 470 117 470 120 7 g
rlabel metal1 470 143 470 146 7 p
<< end >>
