* SPICE3 file created from ckt.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 gnd nor_0/b inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in nor_0/b nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd nor_0/b inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in nor_0/b nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1067 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1068 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a gnd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1071 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1072 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op gnd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1074 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1075 gnd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1076 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1078 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1079 gnd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1080 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a gnd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1083 gnd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1084 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b gnd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1086 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1087 gnd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1088 sumffo_0/ffo_0/nand_7/a clk gnd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1090 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1091 gnd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1092 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a gnd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1095 gnd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1096 z1o sumffo_0/ffo_0/nand_7/a gnd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1098 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1099 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1101 sumffo_0/ffo_0/nand_0/b clk gnd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1102 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_0/xor_0/inv_1/op nor_0/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_0/xor_0/inv_1/op nor_0/b gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 gnd nor_0/b sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 sumffo_0/ffo_0/d nor_0/b sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1115 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1116 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a gnd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1119 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1120 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op gnd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1122 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1123 gnd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1124 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1127 gnd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1128 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a gnd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1130 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1131 gnd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1132 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b gnd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1134 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1135 gnd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1136 sumffo_2/ffo_0/nand_7/a clk gnd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1139 gnd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1140 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a gnd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1143 gnd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1144 z3o sumffo_2/ffo_0/nand_7/a gnd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1146 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1147 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 sumffo_2/ffo_0/nand_0/b clk gnd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1153 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1154 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1155 sumffo_2/ffo_0/d ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1156 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1157 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1158 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1163 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1164 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a gnd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1166 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1167 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1168 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op gnd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1170 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1171 gnd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1172 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a gnd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1179 gnd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1180 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b gnd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1183 gnd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1184 sumffo_1/ffo_0/nand_7/a clk gnd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1186 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1187 gnd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1188 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a gnd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1190 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1191 gnd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1192 z2o sumffo_1/ffo_0/nand_7/a gnd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1194 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1195 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 sumffo_1/ffo_0/nand_0/b clk gnd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1211 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1212 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a gnd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1214 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op gnd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1219 gnd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1220 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1223 gnd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1224 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a gnd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1226 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1227 gnd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1228 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b gnd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1230 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1231 gnd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1232 sumffo_3/ffo_0/nand_7/a clk gnd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1235 gnd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1236 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a gnd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1238 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1239 gnd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1240 z4o sumffo_3/ffo_0/nand_7/a gnd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1245 sumffo_3/ffo_0/nand_0/b clk gnd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1246 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1247 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1248 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1249 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1250 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1251 sumffo_3/ffo_0/d ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1252 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1253 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1254 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1259 gnd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1260 ffo_0/nand_3/b ffo_0/nand_1/a gnd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1262 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1263 gnd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1264 ffo_0/nand_1/a ffo_0/inv_0/op gnd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1266 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1267 gnd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1268 ffo_0/nand_3/a ffo_0/d gnd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1270 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1271 gnd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1272 ffo_0/nand_1/b ffo_0/nand_3/a gnd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1274 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1275 gnd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1276 ffo_0/nand_6/a ffo_0/nand_3/b gnd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1278 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1279 gnd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1280 ffo_0/nand_7/a clk gnd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1282 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1283 gnd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1284 ffo_0/qbar ffo_0/nand_6/a gnd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1286 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1287 gnd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1288 couto ffo_0/nand_7/a gnd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffo_0/inv_0/op ffo_0/d gnd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1293 ffo_0/nand_0/b clk gnd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1294 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1295 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1297 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1298 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1299 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1301 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1303 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1305 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1306 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1307 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1309 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1311 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1313 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1314 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1315 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1317 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1318 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1319 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1320 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1321 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1323 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1325 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1327 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1329 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1330 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1331 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipg_0/pggen_0/nand_0/a_13_n26# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 gnd ffipg_0/ffi_0/q cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 cla_0/g0 ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 cla_0/g0 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1337 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1338 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1339 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 gnd ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1341 ffipg_0/k ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1342 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1343 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1344 ffipg_0/pggen_0/xor_0/a_10_n43# ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/ffi_1/q gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 nor_0/a ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1349 ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/ffi_0/q gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 gnd ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1351 nor_0/a ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 ffipg_0/ffi_0/nand_1/a_13_n26# ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/a gnd ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipg_0/ffi_0/nand_0/a_13_n26# ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 gnd clk ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/inv_0/op gnd ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 ffipg_0/ffi_0/nand_1/a clk ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1361 gnd clk ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1362 ffipg_0/ffi_0/nand_3/a y1in gnd ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 ffipg_0/ffi_0/nand_3/a clk ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipg_0/ffi_0/nand_3/a_13_n26# ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 gnd ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/a gnd ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipg_0/ffi_0/nand_4/a_13_n26# ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1369 gnd ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1370 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/nand_3/b gnd ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1371 ffipg_0/ffi_0/nand_6/a ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 ffipg_0/ffi_0/nand_5/a_13_n26# ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1373 gnd ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1374 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/inv_1/op gnd ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1376 ffipg_0/ffi_0/nand_6/a_13_n26# ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1377 gnd ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1378 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/a gnd ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1380 ffipg_0/ffi_0/nand_7/a_13_n26# ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1381 gnd ffipg_0/ffi_0/qbar ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1382 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a gnd ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1384 ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1385 ffipg_0/ffi_0/inv_0/op y1in gnd ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1386 ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1387 ffipg_0/ffi_0/inv_1/op clk gnd ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipg_0/ffi_1/nand_1/a_13_n26# ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a gnd ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipg_0/ffi_1/nand_0/a_13_n26# ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 gnd clk ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/inv_0/op gnd ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipg_0/ffi_1/nand_1/a clk ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 gnd clk ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipg_0/ffi_1/nand_3/a x1in gnd ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipg_0/ffi_1/nand_3/a clk ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipg_0/ffi_1/nand_3/a_13_n26# ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 gnd ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/a gnd ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipg_0/ffi_1/nand_4/a_13_n26# ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 gnd ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_3/b gnd ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipg_0/ffi_1/nand_5/a_13_n26# ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 gnd ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/inv_1/op gnd ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipg_0/ffi_1/nand_6/a_13_n26# ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 gnd ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_6/a gnd ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipg_0/ffi_1/nand_7/a_13_n26# ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1417 gnd ffipg_0/ffi_1/qbar ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1418 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a gnd ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1421 ffipg_0/ffi_1/inv_0/op x1in gnd ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1422 ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1423 ffipg_0/ffi_1/inv_1/op clk gnd ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1425 ffo_0/d inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1426 ffipg_1/pggen_0/nand_0/a_13_n26# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1427 gnd ffipg_1/ffi_0/q cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 cla_0/l ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 cla_0/l ffipg_1/ffi_0/q ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1431 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1433 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1434 gnd ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1435 ffipg_1/k ffipg_1/ffi_0/q ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1436 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1437 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1438 ffipg_1/pggen_0/xor_0/a_10_n43# ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_1/q gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1441 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 cla_1/p0 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1443 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/ffi_0/q gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 gnd ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1445 cla_1/p0 ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 ffipg_1/ffi_0/nand_1/a_13_n26# ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1447 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1448 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a gnd ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1449 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1450 ffipg_1/ffi_0/nand_0/a_13_n26# ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1451 gnd clk ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1452 ffipg_1/ffi_0/nand_1/a ffipg_1/ffi_0/inv_0/op gnd ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 ffipg_1/ffi_0/nand_1/a clk ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1455 gnd clk ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1456 ffipg_1/ffi_0/nand_3/a y2in gnd ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 ffipg_1/ffi_0/nand_3/a clk ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1458 ffipg_1/ffi_0/nand_3/a_13_n26# ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1459 gnd ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1460 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/a gnd ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1461 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 ffipg_1/ffi_0/nand_4/a_13_n26# ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1463 gnd ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1464 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_3/b gnd ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1466 ffipg_1/ffi_0/nand_5/a_13_n26# ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1467 gnd ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1468 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/inv_1/op gnd ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1470 ffipg_1/ffi_0/nand_6/a_13_n26# ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 gnd ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/a gnd ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 ffipg_1/ffi_0/nand_7/a_13_n26# ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 gnd ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/a gnd ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 ffipg_1/ffi_0/q ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1479 ffipg_1/ffi_0/inv_0/op y2in gnd ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1480 ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1481 ffipg_1/ffi_0/inv_1/op clk gnd ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 ffipg_1/ffi_1/nand_1/a_13_n26# ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a gnd ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 ffipg_1/ffi_1/nand_0/a_13_n26# ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 gnd clk ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 ffipg_1/ffi_1/nand_1/a ffipg_1/ffi_1/inv_0/op gnd ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 ffipg_1/ffi_1/nand_1/a clk ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 gnd clk ffipg_1/ffi_1/nand_3/a ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 ffipg_1/ffi_1/nand_3/a x2in gnd ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 ffipg_1/ffi_1/nand_3/a clk ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 ffipg_1/ffi_1/nand_3/a_13_n26# ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 gnd ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/a gnd ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 ffipg_1/ffi_1/nand_4/a_13_n26# ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 gnd ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_3/b gnd ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 ffipg_1/ffi_1/nand_5/a_13_n26# ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1503 gnd ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1504 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/inv_1/op gnd ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1505 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 ffipg_1/ffi_1/nand_6/a_13_n26# ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1507 gnd ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1508 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a gnd ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 ffipg_1/ffi_1/nand_7/a_13_n26# ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1511 gnd ffipg_1/ffi_1/qbar ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1512 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a gnd ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1513 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1514 ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1515 ffipg_1/ffi_1/inv_0/op x2in gnd ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1516 ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1517 ffipg_1/ffi_1/inv_1/op clk gnd ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1518 ffipg_2/pggen_0/nand_0/a_13_n26# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 gnd ffipg_2/ffi_0/q cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1520 cla_0/l ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 cla_0/l ffipg_2/ffi_0/q ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1523 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1524 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1525 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 gnd ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1527 ffipg_2/k ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1528 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1529 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1530 ffipg_2/pggen_0/xor_0/a_10_n43# ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/ffi_1/q gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1534 cla_2/p0 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1535 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/ffi_0/q gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 gnd ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1537 cla_2/p0 ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 ffipg_2/ffi_0/nand_1/a_13_n26# ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a gnd ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 ffipg_2/ffi_0/nand_0/a_13_n26# ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 gnd clk ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/inv_0/op gnd ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 ffipg_2/ffi_0/nand_1/a clk ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 gnd clk ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 ffipg_2/ffi_0/nand_3/a y3in gnd ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 ffipg_2/ffi_0/nand_3/a clk ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 ffipg_2/ffi_0/nand_3/a_13_n26# ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1551 gnd ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1552 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/a gnd ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 ffipg_2/ffi_0/nand_4/a_13_n26# ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1555 gnd ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1556 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_3/b gnd ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 ffipg_2/ffi_0/nand_5/a_13_n26# ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1559 gnd ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1560 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/inv_1/op gnd ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1561 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1562 ffipg_2/ffi_0/nand_6/a_13_n26# ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1563 gnd ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1564 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_6/a gnd ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1566 ffipg_2/ffi_0/nand_7/a_13_n26# ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 gnd ffipg_2/ffi_0/qbar ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 ffipg_2/ffi_0/q ffipg_2/ffi_0/nand_7/a gnd ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1571 ffipg_2/ffi_0/inv_0/op y3in gnd ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1572 ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1573 ffipg_2/ffi_0/inv_1/op clk gnd ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 ffipg_2/ffi_1/nand_1/a_13_n26# ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/a gnd ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 ffipg_2/ffi_1/nand_0/a_13_n26# ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 gnd clk ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/inv_0/op gnd ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 ffipg_2/ffi_1/nand_1/a clk ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 gnd clk ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 ffipg_2/ffi_1/nand_3/a x3in gnd ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 ffipg_2/ffi_1/nand_3/a clk ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 ffipg_2/ffi_1/nand_3/a_13_n26# ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 gnd ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/a gnd ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 ffipg_2/ffi_1/nand_4/a_13_n26# ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 gnd ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_3/b gnd ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 ffipg_2/ffi_1/nand_5/a_13_n26# ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 gnd ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/inv_1/op gnd ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 ffipg_2/ffi_1/nand_6/a_13_n26# ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1599 gnd ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1600 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/a gnd ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1601 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 ffipg_2/ffi_1/nand_7/a_13_n26# ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1603 gnd ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1604 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/a gnd ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1605 ffipg_2/ffi_1/q ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1607 ffipg_2/ffi_1/inv_0/op x3in gnd ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1608 ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1609 ffipg_2/ffi_1/inv_1/op clk gnd ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1610 ffi_0/nand_1/a_13_n26# ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1611 gnd ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1612 ffi_0/nand_3/b ffi_0/nand_1/a gnd ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1614 ffi_0/nand_0/a_13_n26# ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 gnd clk ffi_0/nand_1/a ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 ffi_0/nand_1/a ffi_0/inv_0/op gnd ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 ffi_0/nand_1/a clk ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 gnd clk ffi_0/nand_3/a ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 ffi_0/nand_3/a cinin gnd ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 ffi_0/nand_3/a clk ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 ffi_0/nand_3/a_13_n26# ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 gnd ffi_0/nand_3/b ffi_0/nand_1/b ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 ffi_0/nand_1/b ffi_0/nand_3/a gnd ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 ffi_0/nand_1/b ffi_0/nand_3/b ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 ffi_0/nand_4/a_13_n26# ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 gnd ffi_0/inv_1/op ffi_0/nand_6/a ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 ffi_0/nand_6/a ffi_0/nand_3/b gnd ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 ffi_0/nand_6/a ffi_0/inv_1/op ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 ffi_0/nand_5/a_13_n26# ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 gnd ffi_0/nand_1/b ffi_0/nand_7/a ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 ffi_0/nand_7/a ffi_0/inv_1/op gnd ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 ffi_0/nand_7/a ffi_0/nand_1/b ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 ffi_0/nand_6/a_13_n26# ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 gnd ffi_0/q nor_0/b ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 nor_0/b ffi_0/nand_6/a gnd ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 nor_0/b ffi_0/q ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 ffi_0/nand_7/a_13_n26# ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 gnd nor_0/b ffi_0/q ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 ffi_0/q ffi_0/nand_7/a gnd ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 ffi_0/q nor_0/b ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1643 ffi_0/inv_0/op cinin gnd ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1644 ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1645 ffi_0/inv_1/op clk gnd ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 ffipg_3/pggen_0/nand_0/a_13_n26# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1647 gnd ffipg_3/ffi_0/q cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1648 cla_2/g1 ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1649 cla_2/g1 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 gnd ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 ffipg_3/k ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 ffipg_3/pggen_0/xor_0/a_10_n43# ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/ffi_1/q gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 cla_2/p1 ffipg_3/ffi_1/q ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1663 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/ffi_0/q gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 gnd ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1665 cla_2/p1 ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1666 ffipg_3/ffi_0/nand_1/a_13_n26# ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/a gnd ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffipg_3/ffi_0/nand_0/a_13_n26# ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 gnd clk ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/inv_0/op gnd ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffipg_3/ffi_0/nand_1/a clk ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 gnd clk ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffipg_3/ffi_0/nand_3/a y4in gnd ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffipg_3/ffi_0/nand_3/a clk ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffipg_3/ffi_0/nand_3/a_13_n26# ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 gnd ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/a gnd ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffipg_3/ffi_0/nand_4/a_13_n26# ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 gnd ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_3/b gnd ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffipg_3/ffi_0/nand_5/a_13_n26# ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 gnd ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/inv_1/op gnd ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffipg_3/ffi_0/nand_6/a_13_n26# ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 gnd ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/a gnd ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffipg_3/ffi_0/nand_7/a_13_n26# ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1695 gnd ffipg_3/ffi_0/qbar ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1696 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_7/a gnd ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1697 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 ffipg_3/ffi_0/inv_0/op y4in gnd ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 ffipg_3/ffi_0/inv_1/op clk gnd ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 ffipg_3/ffi_1/nand_1/a_13_n26# ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1703 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1704 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/a gnd ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1705 ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1706 ffipg_3/ffi_1/nand_0/a_13_n26# ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1707 gnd clk ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1708 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/inv_0/op gnd ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1709 ffipg_3/ffi_1/nand_1/a clk ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1711 gnd clk ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1712 ffipg_3/ffi_1/nand_3/a x4in gnd ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1713 ffipg_3/ffi_1/nand_3/a clk ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1714 ffipg_3/ffi_1/nand_3/a_13_n26# ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1715 gnd ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1716 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/a gnd ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1717 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1718 ffipg_3/ffi_1/nand_4/a_13_n26# ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1719 gnd ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1720 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_3/b gnd ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1721 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 ffipg_3/ffi_1/nand_5/a_13_n26# ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1723 gnd ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1724 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/inv_1/op gnd ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1725 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1726 ffipg_3/ffi_1/nand_6/a_13_n26# ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1727 gnd ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1728 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/a gnd ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1730 ffipg_3/ffi_1/nand_7/a_13_n26# ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1731 gnd ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1732 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/a gnd ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 ffipg_3/ffi_1/q ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 ffipg_3/ffi_1/inv_0/op x4in gnd ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffipg_3/ffi_1/inv_1/op clk gnd ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 ffipg_0/ffi_1/inv_1/w_0_6# gnd 0.06fF
C1 gnd ffipg_3/ffi_1/nand_5/w_0_0# 0.10fF
C2 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C3 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# 0.04fF
C4 gnd ffo_0/nand_1/b 0.57fF
C5 gnd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C6 sumffo_1/ffo_0/d sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C7 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_1/w_0_6# 0.03fF
C8 inv_5/in gnd 0.49fF
C9 cla_1/l nand_2/b 0.31fF
C10 gnd inv_1/in 0.33fF
C11 ffipg_1/ffi_1/q ffipg_1/ffi_1/qbar 0.32fF
C12 ffipg_1/pggen_0/nand_0/w_0_0# ffipg_1/ffi_0/q 0.06fF
C13 clk ffo_0/nand_0/b 0.04fF
C14 sumffo_2/ffo_0/nand_0/b clk 0.04fF
C15 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C16 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C17 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C18 nor_0/a cla_0/nor_0/w_0_0# 0.06fF
C19 ffipg_0/ffi_0/nand_5/w_0_0# gnd 0.10fF
C20 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C21 ffipg_0/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C22 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/b 0.32fF
C23 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C24 ffipg_1/ffi_1/nand_3/b gnd 0.74fF
C25 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/d 0.40fF
C26 inv_8/w_0_6# inv_8/in 0.10fF
C27 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_1/q 0.27fF
C28 clk ffipg_1/ffi_1/inv_1/op 0.07fF
C29 y2in ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C30 inv_5/in nor_3/b 0.04fF
C31 sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# 0.02fF
C32 inv_7/op nor_0/b 0.31fF
C33 cla_0/n cla_0/l 0.25fF
C34 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_3/b 0.00fF
C35 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_1/b 0.45fF
C36 ffipg_1/ffi_1/q ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C37 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/k 0.02fF
C38 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C39 ffipg_1/ffi_0/inv_0/w_0_6# ffipg_1/ffi_0/inv_0/op 0.03fF
C40 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/b 0.31fF
C41 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/k 0.21fF
C42 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_6/a 0.31fF
C43 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C44 sumffo_0/ffo_0/nand_4/w_0_0# gnd 0.10fF
C45 cla_0/n gnd 1.20fF
C46 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C47 gnd ffipg_3/ffi_0/nand_3/b 0.74fF
C48 gnd ffipg_1/ffi_1/nand_1/a 0.44fF
C49 sumffo_3/sbar z4o 0.32fF
C50 sumffo_0/xor_0/w_n3_4# gnd 0.12fF
C51 sumffo_0/xor_0/a_10_10# gnd 0.93fF
C52 ffipg_1/ffi_0/inv_0/w_0_6# gnd 0.06fF
C53 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C54 ffipg_0/ffi_1/inv_0/op gnd 0.27fF
C55 gnd sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C56 sumffo_2/ffo_0/nand_1/b clk 0.45fF
C57 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/a 0.06fF
C58 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a 0.31fF
C59 ffipg_0/ffi_0/nand_6/w_0_0# ffipg_0/ffi_0/nand_6/a 0.06fF
C60 ffipg_3/ffi_0/inv_1/op gnd 1.85fF
C61 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_1/b 0.06fF
C62 ffipg_0/k sumffo_0/xor_0/w_n3_4# 0.06fF
C63 sumffo_0/ffo_0/nand_7/a sumffo_0/sbar 0.31fF
C64 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C65 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/inv_1/op 0.13fF
C66 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C67 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op 0.06fF
C68 gnd ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C69 nor_4/b gnd 0.25fF
C70 ffo_0/nand_4/w_0_0# gnd 0.10fF
C71 sumffo_2/sbar gnd 0.62fF
C72 ffipg_1/pggen_0/nor_0/w_0_0# gnd 0.11fF
C73 nor_0/b sumffo_2/xor_0/inv_1/op 0.04fF
C74 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C75 nor_0/b ffi_0/nand_7/a 0.31fF
C76 ffipg_1/ffi_1/inv_1/w_0_6# ffipg_1/ffi_1/inv_1/op 0.04fF
C77 ffipg_0/ffi_0/nand_3/a gnd 0.33fF
C78 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a 0.00fF
C79 sumffo_2/ffo_0/nand_7/w_0_0# z3o 0.04fF
C80 gnd cla_2/n 0.60fF
C81 ffo_0/nand_3/a ffo_0/nand_3/w_0_0# 0.06fF
C82 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C83 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/q 0.04fF
C84 ffipg_2/ffi_1/inv_1/op clk 0.07fF
C85 ffipg_3/ffi_0/nand_1/w_0_0# gnd 0.10fF
C86 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C87 gnd ffipg_0/ffi_0/nand_3/b 0.74fF
C88 ffi_0/q ffi_0/nand_7/w_0_0# 0.04fF
C89 inv_8/in nor_4/a 0.04fF
C90 gnd ffo_0/nand_3/b 0.74fF
C91 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_0/op 0.32fF
C92 gnd sumffo_3/ffo_0/nand_1/a 0.33fF
C93 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C94 cla_2/l cla_0/l 0.37fF
C95 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_1/b 0.31fF
C96 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C97 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/nand_1/b 0.13fF
C98 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op 0.06fF
C99 nor_3/b cla_2/n 0.41fF
C100 ffipg_1/ffi_1/nand_2/w_0_0# clk 0.06fF
C101 gnd ffipg_3/ffi_1/qbar 0.67fF
C102 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.32fF
C103 ffo_0/d ffo_0/inv_0/op 0.04fF
C104 cla_2/l gnd 0.61fF
C105 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# 0.04fF
C106 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_1/b 0.45fF
C107 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a 0.13fF
C108 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b 0.32fF
C109 sumffo_3/xor_0/a_10_10# nor_0/b 0.04fF
C110 clk ffipg_1/ffi_1/nand_0/w_0_0# 0.06fF
C111 ffipg_2/ffi_0/q ffipg_2/ffi_0/qbar 0.32fF
C112 ffipg_1/ffi_0/nand_3/a clk 0.13fF
C113 ffipg_0/ffi_0/inv_1/op ffipg_0/ffi_0/nand_6/a 0.13fF
C114 gnd ffo_0/nand_1/a 0.33fF
C115 sumffo_0/ffo_0/inv_1/w_0_6# sumffo_0/ffo_0/nand_0/b 0.03fF
C116 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C117 cla_2/l nor_3/b 0.10fF
C118 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C119 ffipg_0/ffi_1/q ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C120 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_1/b 0.06fF
C121 ffo_0/nand_6/a ffo_0/nand_6/w_0_0# 0.06fF
C122 sumffo_2/ffo_0/d nor_0/b 0.27fF
C123 ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C124 gnd ffo_0/nand_7/w_0_0# 0.10fF
C125 cla_0/n inv_3/w_0_6# 0.16fF
C126 ffipg_0/ffi_0/nand_7/w_0_0# ffipg_0/ffi_0/nand_7/a 0.06fF
C127 gnd ffipg_3/ffi_0/nand_6/a 0.37fF
C128 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a 0.31fF
C129 sumffo_0/ffo_0/nand_7/a gnd 0.33fF
C130 cla_2/inv_0/op gnd 0.27fF
C131 gnd ffi_0/nand_5/w_0_0# 0.10fF
C132 gnd ffipg_3/ffi_0/q 3.00fF
C133 gnd ffipg_2/ffi_0/nand_2/w_0_0# 0.10fF
C134 sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# 0.02fF
C135 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C136 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C137 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C138 inv_7/op gnd 0.27fF
C139 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C140 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C141 gnd ffo_0/nand_0/w_0_0# 0.10fF
C142 sumffo_0/ffo_0/nand_1/b gnd 0.57fF
C143 ffipg_3/ffi_0/nand_7/w_0_0# gnd 0.10fF
C144 x2in ffipg_1/ffi_1/inv_0/op 0.04fF
C145 ffipg_0/ffi_0/nand_0/w_0_0# gnd 0.10fF
C146 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C147 gnd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C148 ffi_0/inv_1/op ffi_0/nand_1/b 0.45fF
C149 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_1/inv_1/op 0.75fF
C150 nor_0/b sumffo_3/ffo_0/d 0.16fF
C151 clk ffipg_2/ffi_0/nand_1/a 0.13fF
C152 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C153 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C154 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_3/w_0_0# 0.04fF
C155 ffipg_1/ffi_0/nand_3/b gnd 0.74fF
C156 gnd sumffo_2/ffo_0/nand_3/w_0_0# 0.11fF
C157 gnd ffipg_2/ffi_0/nand_1/b 0.57fF
C158 gnd ffipg_3/ffi_1/nand_3/b 0.74fF
C159 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_7/w_0_0# 0.04fF
C160 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C161 cla_2/nor_1/w_0_0# gnd 0.31fF
C162 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C163 cla_1/p0 ffipg_1/k 0.05fF
C164 nor_4/a nor_4/w_0_0# 0.07fF
C165 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C166 ffo_0/nand_6/a gnd 0.33fF
C167 gnd sumffo_2/ffo_0/nand_4/w_0_0# 0.10fF
C168 ffipg_3/ffi_1/inv_0/op x4in 0.04fF
C169 ffipg_1/ffi_1/q ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C170 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C171 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C172 nor_4/b inv_9/in 0.16fF
C173 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C174 sumffo_2/ffo_0/nand_5/w_0_0# clk 0.06fF
C175 clk sumffo_0/ffo_0/nand_3/b 0.33fF
C176 cla_0/l cla_2/g1 0.26fF
C177 nor_0/b sumffo_1/xor_0/w_n3_4# 0.00fF
C178 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/q 0.00fF
C179 x3in clk 0.68fF
C180 ffipg_1/ffi_1/nand_3/w_0_0# gnd 0.11fF
C181 cla_0/g0 cla_1/p0 0.38fF
C182 gnd ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C183 gnd ffi_0/nand_7/a 0.33fF
C184 gnd sumffo_2/xor_0/inv_1/op 0.35fF
C185 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_6/a 0.13fF
C186 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/b 0.32fF
C187 cla_2/g1 gnd 0.65fF
C188 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C189 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C190 sumffo_0/ffo_0/nand_5/w_0_0# clk 0.06fF
C191 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C192 sumffo_0/ffo_0/nand_6/a clk 0.13fF
C193 cla_0/l cla_1/p0 0.09fF
C194 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_3/b 0.06fF
C195 cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C196 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/b 0.32fF
C197 ffipg_0/ffi_0/nand_2/w_0_0# gnd 0.10fF
C198 sumffo_3/xor_0/inv_1/op inv_4/op 0.06fF
C199 ffipg_3/k sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C200 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C201 cla_1/p0 gnd 1.06fF
C202 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_3/b 0.06fF
C203 ffi_0/nand_1/w_0_0# ffi_0/nand_3/b 0.04fF
C204 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C205 gnd ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C206 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C207 sumffo_3/xor_0/a_10_10# gnd 0.93fF
C208 sumffo_1/ffo_0/nand_1/w_0_0# gnd 0.10fF
C209 ffipg_3/ffi_1/nand_3/a ffipg_3/ffi_1/nand_3/b 0.31fF
C210 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C211 inv_3/in nand_2/b 0.13fF
C212 ffi_0/inv_0/op ffi_0/inv_0/w_0_6# 0.03fF
C213 clk ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C214 clk ffipg_1/ffi_0/inv_0/op 0.32fF
C215 ffipg_0/ffi_1/nand_7/w_0_0# gnd 0.10fF
C216 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C217 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C218 y4in ffipg_3/ffi_0/inv_0/op 0.04fF
C219 gnd sumffo_2/ffo_0/inv_1/w_0_6# 0.07fF
C220 gnd ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C221 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C222 clk sumffo_3/ffo_0/nand_6/a 0.13fF
C223 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C224 clk gnd 24.51fF
C225 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/b 0.31fF
C226 ffipg_2/k cla_2/p0 0.05fF
C227 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_4/w_0_0# 0.04fF
C228 inv_1/op inv_1/in 0.04fF
C229 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C230 ffipg_2/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C231 ffi_0/nand_6/w_0_0# gnd 0.10fF
C232 sumffo_2/ffo_0/d gnd 0.41fF
C233 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_5/w_0_0# 0.04fF
C234 ffipg_1/ffi_1/nand_7/a gnd 0.37fF
C235 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/a 0.06fF
C236 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C237 nor_0/b sumffo_1/xor_0/inv_0/op 0.06fF
C238 clk ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C239 nor_2/w_0_0# inv_4/in 0.11fF
C240 sumffo_3/xor_0/inv_1/op ffipg_3/k 0.22fF
C241 ffo_0/inv_0/w_0_6# ffo_0/d 0.06fF
C242 sumffo_0/ffo_0/nand_3/w_0_0# gnd 0.11fF
C243 cla_2/p0 ffipg_2/ffi_0/q 0.03fF
C244 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/qbar 0.00fF
C245 y1in ffipg_0/ffi_0/inv_1/op 0.01fF
C246 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C247 sumffo_1/xor_0/w_n3_4# ffipg_1/k 0.06fF
C248 ffipg_2/ffi_0/inv_0/w_0_6# y3in 0.06fF
C249 clk ffi_0/inv_1/w_0_6# 0.06fF
C250 sumffo_0/ffo_0/nand_0/a_13_n26# gnd 0.01fF
C251 x1in ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C252 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/ffi_1/q 0.06fF
C253 gnd sumffo_3/ffo_0/d 0.41fF
C254 ffipg_2/k nand_2/b 0.06fF
C255 cinin clk 0.68fF
C256 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C257 ffipg_1/ffi_1/q ffipg_1/ffi_0/q 0.73fF
C258 clk ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C259 nor_0/w_0_0# nor_0/b 0.23fF
C260 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C261 sumffo_1/ffo_0/nand_6/a clk 0.13fF
C262 gnd sumffo_1/ffo_0/nand_2/w_0_0# 0.10fF
C263 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_3/b 0.00fF
C264 ffi_0/nand_1/w_0_0# gnd 0.10fF
C265 ffipg_1/ffi_1/inv_1/w_0_6# gnd 0.06fF
C266 sumffo_0/ffo_0/nand_3/a gnd 0.33fF
C267 ffipg_3/ffi_1/nand_3/a clk 0.13fF
C268 cla_2/p1 ffipg_3/k 0.05fF
C269 ffipg_2/ffi_1/q ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C270 sumffo_3/sbar sumffo_3/ffo_0/nand_7/a 0.31fF
C271 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_1/b 0.45fF
C272 sumffo_2/ffo_0/nand_6/w_0_0# gnd 0.10fF
C273 ffipg_3/k ffipg_3/ffi_1/q 0.46fF
C274 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/w_0_0# 0.04fF
C275 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_3/b 0.04fF
C276 ffipg_3/ffi_0/nand_1/b ffipg_3/ffi_0/nand_5/w_0_0# 0.06fF
C277 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/w_0_0# 0.04fF
C278 couto ffo_0/nand_7/w_0_0# 0.04fF
C279 gnd sumffo_1/xor_0/w_n3_4# 0.12fF
C280 ffipg_2/k ffipg_2/ffi_0/q 0.07fF
C281 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/a 0.00fF
C282 nand_2/b inv_2/w_0_6# 0.03fF
C283 gnd ffipg_3/ffi_0/nand_2/w_0_0# 0.10fF
C284 ffipg_3/ffi_0/nand_0/w_0_0# ffipg_3/ffi_0/inv_0/op 0.06fF
C285 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/b 0.31fF
C286 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/a 0.06fF
C287 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/ffi_0/q 0.06fF
C288 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/w_0_0# 0.04fF
C289 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C290 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C291 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/w_0_0# 0.06fF
C292 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C293 sumffo_2/ffo_0/nand_1/a gnd 0.33fF
C294 ffipg_2/ffi_1/nand_3/b ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C295 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_6/w_0_0# 0.06fF
C296 gnd sumffo_3/ffo_0/nand_6/w_0_0# 0.10fF
C297 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C298 cla_2/nand_0/a_13_n26# gnd 0.01fF
C299 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_3/b 0.00fF
C300 gnd ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C301 gnd ffipg_0/ffi_1/nand_1/b 0.57fF
C302 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C303 cla_0/l cla_0/nand_0/w_0_0# 0.06fF
C304 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_1/b 0.13fF
C305 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/qbar 0.04fF
C306 sumffo_1/ffo_0/d nor_0/b 0.27fF
C307 sumffo_0/ffo_0/d clk 0.25fF
C308 ffipg_1/ffi_0/inv_1/op ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C309 ffipg_0/ffi_0/q ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C310 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/a 0.00fF
C311 gnd ffipg_3/ffi_1/inv_1/op 1.85fF
C312 gnd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C313 cla_0/nand_0/w_0_0# gnd 0.10fF
C314 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/ffi_1/q 0.06fF
C315 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/b 0.31fF
C316 gnd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C317 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C318 inv_5/in inv_5/w_0_6# 0.10fF
C319 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C320 ffo_0/nand_1/w_0_0# ffo_0/nand_1/a 0.06fF
C321 ffipg_2/ffi_0/inv_0/w_0_6# ffipg_2/ffi_0/inv_0/op 0.03fF
C322 ffipg_0/ffi_0/q cla_0/g0 0.13fF
C323 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C324 couto ffo_0/nand_6/a 0.31fF
C325 sumffo_0/ffo_0/inv_0/op gnd 0.27fF
C326 ffipg_3/ffi_0/inv_0/w_0_6# gnd 0.06fF
C327 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C328 ffipg_0/ffi_0/inv_0/op gnd 0.27fF
C329 gnd sumffo_3/ffo_0/nand_3/a 0.33fF
C330 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C331 ffipg_3/ffi_0/inv_1/w_0_6# gnd 0.06fF
C332 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k 0.52fF
C333 gnd ffipg_1/ffi_0/inv_1/op 1.85fF
C334 sumffo_1/xor_0/inv_0/op gnd 0.32fF
C335 ffipg_0/ffi_0/q gnd 3.00fF
C336 cla_0/n inv_5/w_0_6# 0.06fF
C337 nor_0/w_0_0# cla_0/g0 0.06fF
C338 ffipg_1/ffi_0/q ffipg_1/ffi_0/nand_7/w_0_0# 0.04fF
C339 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_5/w_0_0# 0.04fF
C340 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/a 0.06fF
C341 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C342 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C343 ffipg_1/ffi_0/nand_0/w_0_0# ffipg_1/ffi_0/inv_0/op 0.06fF
C344 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_7/w_0_0# 0.06fF
C345 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/ffi_0/q 0.22fF
C346 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C347 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# 0.04fF
C348 ffipg_0/ffi_0/q ffipg_0/k 0.07fF
C349 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_6/a 0.04fF
C350 sumffo_3/ffo_0/nand_4/w_0_0# gnd 0.10fF
C351 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C352 ffipg_1/ffi_0/nand_0/w_0_0# gnd 0.10fF
C353 inv_8/w_0_6# nor_4/a 0.03fF
C354 nor_0/w_0_0# gnd 0.46fF
C355 ffipg_2/ffi_0/nand_1/w_0_0# gnd 0.10fF
C356 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C357 clk ffipg_3/ffi_1/nand_1/a 0.13fF
C358 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/ffi_0/q 0.23fF
C359 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/inv_1/w_0_6# 0.04fF
C360 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/qbar 0.31fF
C361 clk sumffo_1/ffo_0/nand_0/b 0.04fF
C362 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C363 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C364 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k 0.06fF
C365 ffipg_0/ffi_1/nand_0/w_0_0# ffipg_0/ffi_1/inv_0/op 0.06fF
C366 ffipg_2/ffi_0/nand_3/b gnd 0.74fF
C367 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/inv_1/op 0.45fF
C368 cla_0/n cla_1/inv_0/w_0_6# 0.26fF
C369 ffi_0/nand_0/a_13_n26# gnd 0.01fF
C370 gnd ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C371 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/inv_1/op 0.13fF
C372 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C373 ffipg_1/ffi_0/nand_6/a gnd 0.37fF
C374 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C375 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C376 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C377 cla_2/l cla_2/p1 0.02fF
C378 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/inv_1/op 0.33fF
C379 cla_0/n cla_1/l 0.07fF
C380 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# 0.04fF
C381 ffipg_2/k ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C382 gnd sumffo_1/ffo_0/nand_3/b 0.74fF
C383 cla_2/l inv_5/w_0_6# 0.08fF
C384 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/q 0.32fF
C385 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/ffi_1/q 0.27fF
C386 inv_2/in nand_2/b 0.34fF
C387 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_5/w_0_0# 0.04fF
C388 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/d 0.06fF
C389 sumffo_2/ffo_0/inv_0/w_0_6# gnd 0.07fF
C390 ffipg_3/ffi_1/nand_2/w_0_0# clk 0.06fF
C391 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/ffi_0/q 0.20fF
C392 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C393 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C394 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C395 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_0/q 0.22fF
C396 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_6/a 0.04fF
C397 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C398 ffipg_0/ffi_1/nand_1/b ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C399 ffipg_2/pggen_0/xor_0/a_10_10# gnd 0.93fF
C400 gnd sumffo_1/ffo_0/nand_7/a 0.33fF
C401 ffipg_2/ffi_1/nand_1/b gnd 0.57fF
C402 sumffo_3/ffo_0/inv_1/w_0_6# gnd 0.06fF
C403 sumffo_1/ffo_0/d gnd 0.41fF
C404 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/op 0.04fF
C405 gnd nor_1/b 0.35fF
C406 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C407 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/b 0.06fF
C408 ffo_0/nand_5/w_0_0# clk 0.06fF
C409 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C410 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C411 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C412 gnd z3o 0.80fF
C413 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C414 cla_1/nor_0/w_0_0# gnd 0.31fF
C415 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/ffi_1/q 0.06fF
C416 ffipg_2/ffi_0/nand_3/a ffipg_2/ffi_0/nand_2/w_0_0# 0.04fF
C417 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/q 0.32fF
C418 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C419 cla_2/inv_0/in cla_2/g1 0.04fF
C420 cla_0/inv_0/op cla_0/nand_0/w_0_0# 0.06fF
C421 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/qbar 0.04fF
C422 cla_2/p1 ffipg_3/ffi_0/q 0.03fF
C423 ffipg_0/ffi_1/nand_3/a clk 0.13fF
C424 ffipg_2/ffi_1/nand_1/w_0_0# gnd 0.10fF
C425 x1in gnd 0.22fF
C426 inv_2/in inv_2/w_0_6# 0.10fF
C427 ffipg_3/ffi_0/nand_1/a clk 0.13fF
C428 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C429 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/nand_7/a 0.06fF
C430 nor_0/w_0_0# inv_0/in 0.11fF
C431 ffipg_3/ffi_0/q ffipg_3/ffi_1/q 0.73fF
C432 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C433 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/sbar 0.04fF
C434 sumffo_2/ffo_0/nand_3/b clk 0.33fF
C435 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C436 cla_0/nand_0/a_13_n26# gnd 0.00fF
C437 gnd ffipg_3/ffi_1/nand_1/b 0.57fF
C438 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/ffi_1/q 0.06fF
C439 ffi_0/nand_6/w_0_0# ffi_0/nand_6/a 0.06fF
C440 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C441 inv_4/in inv_4/op 0.04fF
C442 ffo_0/nand_6/a ffo_0/qbar 0.00fF
C443 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C444 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C445 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_1/op 0.08fF
C446 ffipg_2/ffi_1/q ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C447 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C448 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C449 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/inv_0/op 0.08fF
C450 gnd ffo_0/nand_0/b 0.58fF
C451 sumffo_2/ffo_0/nand_0/b gnd 0.63fF
C452 ffipg_3/ffi_1/inv_0/op ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C453 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C454 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C455 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C456 ffipg_3/ffi_0/nand_3/a clk 0.13fF
C457 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/ffo_0/nand_6/a 0.06fF
C458 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C459 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C460 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C461 gnd ffipg_1/ffi_1/inv_1/op 1.85fF
C462 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C463 x1in ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C464 sumffo_0/ffo_0/nand_0/w_0_0# gnd 0.10fF
C465 cla_2/p1 cla_2/g1 0.00fF
C466 ffipg_0/ffi_0/nand_7/a ffipg_0/ffi_0/qbar 0.31fF
C467 ffipg_2/ffi_1/inv_1/op x3in 0.01fF
C468 y2in ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C469 ffipg_0/ffi_1/nand_1/a clk 0.13fF
C470 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C471 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_1/b 0.04fF
C472 ffipg_0/ffi_1/inv_0/w_0_6# gnd 0.06fF
C473 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C474 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C475 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a 0.31fF
C476 cla_0/l inv_7/w_0_6# 0.06fF
C477 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_1/b 0.04fF
C478 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C479 nor_4/b nor_4/w_0_0# 0.06fF
C480 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_3/b 0.04fF
C481 gnd ffipg_3/ffi_1/nand_6/w_0_0# 0.10fF
C482 sumffo_2/ffo_0/nand_1/b gnd 0.57fF
C483 inv_7/w_0_6# gnd 0.15fF
C484 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_3/a 0.31fF
C485 gnd ffipg_1/ffi_0/nand_4/w_0_0# 0.10fF
C486 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C487 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_0/q 0.22fF
C488 clk ffipg_2/ffi_1/inv_0/op 0.32fF
C489 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/sbar 0.04fF
C490 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/inv_1/op 0.06fF
C491 ffipg_2/ffi_0/nand_6/w_0_0# ffipg_2/ffi_0/q 0.06fF
C492 clk ffipg_2/ffi_0/nand_3/a 0.13fF
C493 sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d 0.52fF
C494 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k 0.06fF
C495 gnd ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C496 ffipg_3/ffi_1/nand_7/a gnd 0.37fF
C497 gnd ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C498 nor_0/b ffipg_1/k 0.06fF
C499 clk ffipg_3/ffi_0/inv_0/op 0.32fF
C500 ffipg_2/ffi_1/inv_1/op gnd 1.85fF
C501 ffipg_2/ffi_1/nand_3/a clk 0.13fF
C502 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a 0.00fF
C503 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C504 cla_2/nand_0/w_0_0# gnd 0.18fF
C505 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C506 clk x4in 0.68fF
C507 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/ffi_0/q 0.12fF
C508 clk ffipg_0/ffi_0/inv_1/op 0.07fF
C509 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C510 ffipg_1/ffi_0/nand_6/w_0_0# gnd 0.10fF
C511 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C512 cla_2/p0 ffipg_3/k 0.06fF
C513 ffipg_3/ffi_0/nand_3/a ffipg_3/ffi_0/nand_2/w_0_0# 0.04fF
C514 sumffo_1/ffo_0/nand_7/a sumffo_1/sbar 0.31fF
C515 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C516 sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d 0.06fF
C517 sumffo_0/ffo_0/inv_1/w_0_6# clk 0.06fF
C518 sumffo_0/ffo_0/nand_1/w_0_0# gnd 0.10fF
C519 cla_0/nor_1/w_0_0# cla_0/l 0.02fF
C520 cla_0/g0 nor_0/b 0.08fF
C521 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_6/w_0_0# 0.06fF
C522 ffipg_1/ffi_1/nand_2/w_0_0# gnd 0.10fF
C523 cla_0/nor_1/w_0_0# gnd 0.31fF
C524 gnd ffipg_1/ffi_1/nand_0/w_0_0# 0.10fF
C525 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/ffo_0/nand_7/a 0.06fF
C526 ffipg_1/ffi_0/nand_3/a gnd 0.33fF
C527 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C528 nor_1/w_0_0# inv_1/in 0.11fF
C529 ffi_0/nand_5/w_0_0# ffi_0/nand_1/b 0.06fF
C530 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_1/b 0.04fF
C531 ffipg_0/ffi_1/nand_0/w_0_0# clk 0.06fF
C532 cla_1/p0 cla_1/l 0.16fF
C533 cla_0/l nor_0/b 0.33fF
C534 clk ffi_0/nand_0/w_0_0# 0.06fF
C535 ffipg_1/pggen_0/xor_0/inv_0/op gnd 0.32fF
C536 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C537 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_1/w_0_6# 0.03fF
C538 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a 0.00fF
C539 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# 0.04fF
C540 nor_0/b gnd 2.12fF
C541 ffi_0/nand_3/a clk 0.13fF
C542 ffipg_1/pggen_0/nand_0/w_0_0# cla_1/p0 0.24fF
C543 sumffo_0/ffo_0/nand_6/a sumffo_0/sbar 0.00fF
C544 nor_0/a ffipg_0/pggen_0/nand_0/w_0_0# 0.24fF
C545 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/b 0.31fF
C546 ffipg_2/ffi_1/inv_1/w_0_6# clk 0.06fF
C547 gnd sumffo_3/ffo_0/nand_0/w_0_0# 0.10fF
C548 sumffo_1/ffo_0/d sumffo_1/ffo_0/nand_0/b 0.40fF
C549 sumffo_0/ffo_0/nand_6/w_0_0# gnd 0.10fF
C550 ffipg_3/ffi_1/nand_1/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C551 nor_1/w_0_0# cla_0/n 0.06fF
C552 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C553 ffipg_0/k nor_0/b 0.19fF
C554 sumffo_0/ffo_0/nand_7/a z1o 0.00fF
C555 ffipg_1/ffi_1/nand_7/a ffipg_1/ffi_1/qbar 0.31fF
C556 ffipg_0/ffi_0/q ffipg_0/ffi_1/q 0.73fF
C557 gnd ffipg_1/ffi_1/nand_6/a 0.37fF
C558 ffipg_1/ffi_1/inv_0/w_0_6# gnd 0.06fF
C559 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C560 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/inv_0/w_0_6# 0.03fF
C561 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# 0.16fF
C562 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/q 0.00fF
C563 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C564 ffo_0/nand_7/a ffo_0/nand_1/b 0.13fF
C565 gnd ffipg_2/ffi_0/nand_1/a 0.44fF
C566 sumffo_2/ffo_0/nand_1/w_0_0# gnd 0.10fF
C567 sumffo_0/sbar gnd 0.62fF
C568 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_1/b 0.31fF
C569 ffi_0/nand_7/a ffi_0/nand_1/b 0.13fF
C570 ffipg_2/ffi_0/nand_5/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C571 gnd ffi_0/nand_3/b 0.74fF
C572 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_6/a 0.13fF
C573 ffipg_0/ffi_1/inv_1/op clk 0.07fF
C574 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_1/b 0.06fF
C575 nor_2/w_0_0# inv_4/op 0.03fF
C576 ffipg_1/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C577 ffi_0/nand_4/w_0_0# ffi_0/nand_3/b 0.06fF
C578 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C579 gnd ffipg_3/ffi_1/nand_7/w_0_0# 0.10fF
C580 ffi_0/q ffi_0/nand_7/a 0.00fF
C581 ffipg_0/ffi_1/nand_6/w_0_0# gnd 0.10fF
C582 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C583 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C584 cla_0/g0 ffipg_1/k 0.06fF
C585 ffo_0/inv_1/w_0_6# clk 0.06fF
C586 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C587 x3in ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C588 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_1/b 0.04fF
C589 clk ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C590 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/nand_7/a 0.06fF
C591 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C592 gnd ffo_0/nand_6/w_0_0# 0.10fF
C593 gnd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C594 sumffo_2/ffo_0/nand_5/w_0_0# gnd 0.10fF
C595 sumffo_0/ffo_0/nand_3/b gnd 0.74fF
C596 ffipg_3/ffi_1/inv_1/op x4in 0.01fF
C597 x3in gnd 0.22fF
C598 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_5/w_0_0# 0.04fF
C599 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C600 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_3/b 0.04fF
C601 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C602 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C603 ffipg_0/pggen_0/nor_0/w_0_0# gnd 0.11fF
C604 gnd ffipg_1/k 0.70fF
C605 sumffo_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C606 sumffo_0/ffo_0/nand_5/w_0_0# gnd 0.10fF
C607 ffipg_3/ffi_0/inv_0/w_0_6# ffipg_3/ffi_0/inv_0/op 0.03fF
C608 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/sbar 0.06fF
C609 sumffo_0/ffo_0/nand_6/a gnd 0.33fF
C610 gnd ffipg_1/ffi_0/nand_5/w_0_0# 0.10fF
C611 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C612 sumffo_3/ffo_0/nand_1/w_0_0# gnd 0.10fF
C613 cla_0/n nand_2/b 0.06fF
C614 clk ffi_0/nand_1/a 0.13fF
C615 nor_0/b inv_0/in 0.23fF
C616 cla_0/g0 cla_0/l 0.14fF
C617 y3in ffipg_2/ffi_0/inv_1/op 0.01fF
C618 cla_0/n ffipg_2/k 0.06fF
C619 gnd ffipg_3/ffi_0/nand_1/b 0.57fF
C620 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C621 ffipg_0/k ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C622 inv_6/in nor_3/w_0_0# 0.11fF
C623 ffo_0/inv_0/w_0_6# ffo_0/inv_0/op 0.03fF
C624 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C625 sumffo_0/xor_0/inv_0/w_0_6# ffipg_0/k 0.06fF
C626 cla_0/g0 gnd 1.03fF
C627 ffipg_2/pggen_0/nor_0/w_0_0# ffipg_2/ffi_0/q 0.06fF
C628 sumffo_1/ffo_0/nand_5/w_0_0# clk 0.06fF
C629 y2in clk 0.68fF
C630 ffipg_0/ffi_0/inv_1/w_0_6# clk 0.06fF
C631 ffipg_1/ffi_1/nand_3/w_0_0# ffipg_1/ffi_1/nand_3/a 0.06fF
C632 ffipg_0/ffi_1/nand_7/w_0_0# ffipg_0/ffi_1/qbar 0.06fF
C633 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/ffo_0/nand_7/a 0.06fF
C634 gnd ffipg_2/ffi_1/nand_2/w_0_0# 0.10fF
C635 ffipg_1/ffi_0/nand_7/a gnd 0.37fF
C636 gnd ffipg_1/ffi_0/inv_0/op 0.27fF
C637 gnd sumffo_3/ffo_0/nand_3/b 0.74fF
C638 ffi_0/nand_6/w_0_0# ffi_0/q 0.06fF
C639 cla_2/l cla_2/p0 0.16fF
C640 cla_0/l gnd 3.05fF
C641 gnd ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C642 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_3/a 0.04fF
C643 z3o sumffo_2/ffo_0/nand_7/a 0.00fF
C644 nor_0/b sumffo_3/xor_0/a_38_n43# 0.01fF
C645 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C646 clk ffi_0/nand_2/w_0_0# 0.06fF
C647 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/ffi_0/q 0.06fF
C648 sumffo_3/ffo_0/nand_6/a gnd 0.33fF
C649 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/a 0.00fF
C650 ffi_0/nand_4/w_0_0# gnd 0.10fF
C651 gnd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C652 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/nand_6/a 0.06fF
C653 sumffo_3/ffo_0/d sumffo_3/ffo_0/inv_0/op 0.04fF
C654 ffipg_3/ffi_0/nand_6/w_0_0# ffipg_3/ffi_0/q 0.06fF
C655 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/a 0.31fF
C656 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C657 ffipg_0/k gnd 0.68fF
C658 gnd ffipg_2/ffi_1/nand_0/w_0_0# 0.10fF
C659 ffipg_0/ffi_0/nand_3/b ffipg_0/ffi_0/nand_1/a 0.00fF
C660 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/nand_1/b 0.13fF
C661 ffi_0/nand_1/w_0_0# ffi_0/nand_1/a 0.06fF
C662 ffipg_2/ffi_1/qbar gnd 0.67fF
C663 ffipg_1/ffi_1/q ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C664 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_1/b 0.45fF
C665 gnd nor_3/b 0.33fF
C666 ffi_0/nand_1/w_0_0# ffi_0/nand_1/b 0.06fF
C667 clk ffipg_1/ffi_1/inv_0/op 0.32fF
C668 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a 0.31fF
C669 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/op 0.04fF
C670 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_3/b 0.32fF
C671 gnd ffi_0/inv_1/w_0_6# 0.06fF
C672 clk ffipg_1/ffi_1/nand_3/a 0.13fF
C673 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_7/a 0.13fF
C674 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/nand_3/b 0.06fF
C675 ffo_0/nand_1/b ffo_0/nand_3/w_0_0# 0.04fF
C676 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a 0.13fF
C677 sumffo_1/ffo_0/nand_6/w_0_0# z2o 0.06fF
C678 sumffo_0/xor_0/inv_1/w_0_6# nor_0/b 0.23fF
C679 ffipg_3/ffi_1/nand_4/w_0_0# gnd 0.10fF
C680 ffo_0/nand_7/a ffo_0/nand_7/w_0_0# 0.06fF
C681 cinin gnd 0.22fF
C682 sumffo_0/ffo_0/nand_7/w_0_0# gnd 0.10fF
C683 gnd ffipg_0/ffi_1/nand_2/w_0_0# 0.10fF
C684 ffipg_3/ffi_1/nand_3/w_0_0# gnd 0.11fF
C685 ffipg_3/ffi_0/nand_7/a gnd 0.37fF
C686 ffipg_1/ffi_0/nand_1/b gnd 0.57fF
C687 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/b 0.32fF
C688 sumffo_1/ffo_0/nand_6/a gnd 0.33fF
C689 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C690 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/nand_1/b 0.13fF
C691 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_1/a 0.31fF
C692 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_3/b 0.04fF
C693 ffipg_3/ffi_1/nand_3/a gnd 0.33fF
C694 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b 0.32fF
C695 cla_0/l cla_1/n 0.13fF
C696 ffipg_2/ffi_1/nand_1/a clk 0.13fF
C697 ffipg_2/ffi_0/nand_6/a gnd 0.37fF
C698 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C699 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C700 gnd sumffo_2/ffo_0/nand_3/a 0.33fF
C701 gnd cla_1/n 0.51fF
C702 ffipg_1/ffi_0/inv_1/w_0_6# ffipg_1/ffi_0/inv_1/op 0.04fF
C703 cla_0/l cla_1/inv_0/in 0.23fF
C704 ffipg_1/ffi_1/nand_1/w_0_0# ffipg_1/ffi_1/nand_1/a 0.06fF
C705 gnd ffipg_2/ffi_1/nand_6/a 0.37fF
C706 sumffo_2/ffo_0/nand_2/w_0_0# gnd 0.10fF
C707 cla_1/nand_0/a_13_n26# gnd 0.01fF
C708 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C709 gnd inv_0/in 0.30fF
C710 cla_1/inv_0/in gnd 0.34fF
C711 ffipg_0/ffi_0/nand_0/w_0_0# ffipg_0/ffi_0/nand_1/a 0.04fF
C712 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C713 clk ffi_0/inv_0/op 0.32fF
C714 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C715 nor_4/b nor_4/a 0.42fF
C716 sumffo_0/ffo_0/d gnd 0.41fF
C717 gnd inv_3/w_0_6# 0.17fF
C718 ffipg_3/ffi_1/nand_3/w_0_0# ffipg_3/ffi_1/nand_3/a 0.06fF
C719 ffipg_3/pggen_0/nand_0/w_0_0# ffipg_3/ffi_1/q 0.06fF
C720 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/a 0.00fF
C721 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_1/a 0.00fF
C722 clk ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C723 inv_7/op inv_8/w_0_6# 0.06fF
C724 ffipg_2/ffi_0/nand_0/w_0_0# ffipg_2/ffi_0/inv_0/op 0.06fF
C725 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C726 cla_1/p0 cla_2/p0 0.24fF
C727 gnd ffipg_0/ffi_0/nand_1/b 0.57fF
C728 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C729 inv_9/in gnd 0.33fF
C730 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C731 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C732 gnd ffipg_0/ffi_1/nand_1/w_0_0# 0.10fF
C733 y2in ffipg_1/ffi_0/inv_1/op 0.01fF
C734 ffo_0/nand_3/b ffo_0/nand_3/w_0_0# 0.06fF
C735 cla_0/l cla_0/inv_0/op 0.35fF
C736 couto ffo_0/nand_6/w_0_0# 0.06fF
C737 ffo_0/d ffo_0/nand_0/b 0.40fF
C738 ffi_0/nand_7/w_0_0# ffi_0/nand_7/a 0.06fF
C739 ffipg_0/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C740 nor_0/b ffi_0/nand_6/a 0.00fF
C741 ffipg_2/k sumffo_2/xor_0/inv_1/op 0.22fF
C742 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C743 cla_0/inv_0/op gnd 0.27fF
C744 ffipg_2/ffi_0/q ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C745 cla_0/n cla_1/inv_0/op 0.06fF
C746 cla_1/p0 ffipg_1/ffi_0/q 0.03fF
C747 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C748 gnd ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C749 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C750 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C751 ffipg_0/pggen_0/xor_0/inv_1/op gnd 0.35fF
C752 ffo_0/nand_3/a ffo_0/nand_0/b 0.13fF
C753 gnd sumffo_1/sbar 0.62fF
C754 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C755 gnd ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C756 inv_7/op inv_7/in 0.04fF
C757 cla_1/p0 ffipg_2/k 0.06fF
C758 gnd nor_2/b 0.32fF
C759 sumffo_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C760 ffipg_3/ffi_1/nand_6/w_0_0# ffipg_3/ffi_1/q 0.06fF
C761 ffi_0/inv_1/op ffi_0/nand_5/w_0_0# 0.06fF
C762 ffipg_2/ffi_1/nand_3/w_0_0# gnd 0.11fF
C763 ffipg_0/ffi_0/nand_7/w_0_0# gnd 0.10fF
C764 sumffo_2/xor_0/inv_1/w_0_6# gnd 0.06fF
C765 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/nand_3/a 0.04fF
C766 ffipg_1/ffi_1/q cla_1/p0 0.22fF
C767 ffi_0/nand_3/w_0_0# ffi_0/nand_3/b 0.06fF
C768 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k 0.52fF
C769 gnd ffipg_3/ffi_1/nand_1/a 0.44fF
C770 sumffo_3/ffo_0/inv_0/w_0_6# gnd 0.07fF
C771 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C772 ffipg_0/ffi_1/inv_1/op x1in 0.01fF
C773 ffipg_0/ffi_1/nand_6/a ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C774 clk ffipg_0/ffi_0/nand_1/a 0.13fF
C775 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_3/b 0.04fF
C776 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C777 clk ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C778 sumffo_3/xor_0/inv_1/op nor_0/b 0.04fF
C779 y3in ffipg_2/ffi_0/inv_0/op 0.04fF
C780 clk ffipg_1/ffi_0/nand_1/a 0.13fF
C781 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C782 couto gnd 0.80fF
C783 sumffo_1/ffo_0/nand_0/b gnd 0.62fF
C784 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/q 0.00fF
C785 gnd sumffo_1/ffo_0/nand_1/a 0.44fF
C786 ffipg_3/ffi_1/inv_0/w_0_6# x4in 0.06fF
C787 nor_0/b sumffo_2/xor_0/a_10_10# 0.04fF
C788 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C789 ffipg_2/pggen_0/nand_0/w_0_0# ffipg_2/ffi_0/q 0.06fF
C790 clk sumffo_3/ffo_0/nand_0/b 0.04fF
C791 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C792 ffipg_0/ffi_0/q ffipg_0/ffi_0/qbar 0.32fF
C793 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_2/w_0_0# 0.06fF
C794 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/w_n3_4# 0.06fF
C795 sumffo_1/ffo_0/nand_6/a sumffo_1/sbar 0.00fF
C796 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C797 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_7/a 0.04fF
C798 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C799 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C800 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/a 0.00fF
C801 ffipg_1/ffi_1/nand_3/w_0_0# ffipg_1/ffi_1/nand_1/b 0.04fF
C802 clk x2in 0.68fF
C803 ffipg_0/ffi_1/nand_6/w_0_0# ffipg_0/ffi_1/q 0.06fF
C804 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C805 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C806 ffipg_0/ffi_1/nand_3/w_0_0# ffipg_0/ffi_1/nand_1/b 0.04fF
C807 ffipg_3/ffi_1/nand_2/w_0_0# gnd 0.10fF
C808 ffo_0/inv_1/w_0_6# ffo_0/nand_0/b 0.03fF
C809 ffipg_3/k inv_4/op 0.09fF
C810 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C811 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C812 nor_4/b nor_3/w_0_0# 0.03fF
C813 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C814 sumffo_2/ffo_0/nand_6/a gnd 0.33fF
C815 x3in ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C816 nor_3/w_0_0# cla_2/n 0.06fF
C817 ffipg_3/ffi_0/nand_1/a ffipg_3/ffi_0/nand_1/b 0.31fF
C818 ffo_0/nand_5/w_0_0# gnd 0.10fF
C819 gnd ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C820 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C821 ffipg_0/ffi_1/q ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C822 nor_2/b cla_1/n 0.39fF
C823 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/d 0.40fF
C824 sumffo_2/xor_0/inv_0/op nor_0/b 0.06fF
C825 sumffo_2/xor_0/w_n3_4# nor_0/b 0.00fF
C826 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C827 ffipg_2/ffi_1/inv_1/w_0_6# ffipg_2/ffi_1/inv_1/op 0.04fF
C828 ffi_0/nand_3/w_0_0# gnd 0.11fF
C829 ffipg_1/ffi_1/nand_7/w_0_0# gnd 0.10fF
C830 nor_4/b inv_6/in 0.04fF
C831 ffipg_0/ffi_1/nand_3/a gnd 0.33fF
C832 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C833 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_3/b 0.32fF
C834 inv_6/in cla_2/n 0.02fF
C835 gnd ffo_0/nand_1/w_0_0# 0.10fF
C836 ffipg_3/k sumffo_3/xor_0/inv_0/op 0.20fF
C837 inv_1/op gnd 0.58fF
C838 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C839 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C840 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/a 0.06fF
C841 nor_0/a cla_1/p0 0.24fF
C842 ffipg_3/ffi_0/nand_1/a gnd 0.44fF
C843 gnd ffi_0/nand_6/a 0.33fF
C844 ffi_0/nand_4/w_0_0# ffi_0/nand_6/a 0.04fF
C845 nor_2/b inv_3/w_0_6# 0.03fF
C846 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C847 gnd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C848 sumffo_2/ffo_0/nand_3/b gnd 0.74fF
C849 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/inv_1/op 0.13fF
C850 ffipg_2/ffi_0/nand_1/b ffipg_2/ffi_0/inv_1/op 0.45fF
C851 ffi_0/inv_1/op clk 0.93fF
C852 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_7/a 0.13fF
C853 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_0/op 0.08fF
C854 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/nand_7/a 0.13fF
C855 gnd sumffo_2/ffo_0/nand_7/a 0.33fF
C856 ffipg_3/ffi_1/nand_2/w_0_0# ffipg_3/ffi_1/nand_3/a 0.04fF
C857 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# gnd 0.06fF
C858 gnd ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C859 ffipg_2/ffi_1/nand_1/w_0_0# ffipg_2/ffi_1/nand_3/b 0.04fF
C860 ffipg_0/ffi_1/q gnd 2.24fF
C861 ffo_0/qbar ffo_0/nand_6/w_0_0# 0.04fF
C862 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C863 clk nor_4/a 0.03fF
C864 x3in ffipg_2/ffi_1/inv_0/op 0.04fF
C865 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C866 cla_0/l cla_2/inv_0/in 0.16fF
C867 nor_0/b inv_8/in 0.13fF
C868 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_3/a 0.04fF
C869 y4in ffipg_3/ffi_0/inv_1/op 0.01fF
C870 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C871 ffipg_3/ffi_0/nand_3/a gnd 0.33fF
C872 gnd ffipg_2/ffi_1/q 2.24fF
C873 cla_2/inv_0/in gnd 0.34fF
C874 ffipg_3/ffi_1/q ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C875 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_2/w_0_0# 0.04fF
C876 ffipg_0/ffi_1/q ffipg_0/k 0.46fF
C877 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_1/b 0.31fF
C878 sumffo_0/ffo_0/inv_0/w_0_6# gnd 0.06fF
C879 cla_0/inv_0/w_0_6# gnd 0.06fF
C880 ffipg_1/ffi_1/qbar ffipg_1/ffi_1/nand_6/a 0.00fF
C881 ffipg_0/ffi_1/nand_1/a gnd 0.45fF
C882 gnd ffipg_0/ffi_0/nand_6/w_0_0# 0.10fF
C883 sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# 0.02fF
C884 sumffo_3/xor_0/inv_1/op gnd 0.35fF
C885 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/q 0.32fF
C886 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C887 gnd sumffo_2/xor_0/a_10_10# 0.93fF
C888 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C889 ffipg_0/ffi_0/nand_3/w_0_0# gnd 0.11fF
C890 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a 0.13fF
C891 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C892 sumffo_1/ffo_0/inv_0/op gnd 0.27fF
C893 cla_0/nor_0/w_0_0# gnd 0.31fF
C894 ffi_0/nand_3/a ffi_0/nand_3/b 0.31fF
C895 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C896 ffipg_0/ffi_0/nand_5/w_0_0# ffipg_0/ffi_0/nand_7/a 0.04fF
C897 ffipg_2/ffi_1/inv_0/op gnd 0.27fF
C898 gnd ffo_0/qbar 0.62fF
C899 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C900 gnd z4o 0.80fF
C901 nor_1/w_0_0# nor_1/b 0.06fF
C902 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/ffi_1/q 0.06fF
C903 cla_0/n ffipg_3/k 0.06fF
C904 clk ffipg_2/ffi_0/inv_1/op 0.07fF
C905 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/nand_7/a 0.04fF
C906 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a 0.31fF
C907 sumffo_0/ffo_0/nand_0/b clk 0.04fF
C908 cla_0/l cla_2/p1 0.30fF
C909 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C910 ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_2/w_0_0# 0.04fF
C911 gnd ffipg_2/ffi_0/nand_3/a 0.33fF
C912 gnd ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C913 sumffo_0/ffo_0/nand_2/w_0_0# gnd 0.10fF
C914 ffipg_3/ffi_0/nand_3/b ffipg_3/ffi_0/nand_4/w_0_0# 0.06fF
C915 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C916 gnd ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C917 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C918 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C919 cla_2/p1 gnd 1.00fF
C920 nor_0/w_0_0# nand_2/b 0.04fF
C921 ffipg_1/ffi_0/nand_0/w_0_0# ffipg_1/ffi_0/nand_1/a 0.04fF
C922 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_1/op 0.52fF
C923 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C924 ffipg_3/ffi_0/qbar ffipg_3/ffi_0/nand_6/a 0.00fF
C925 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/ffi_1/q 0.06fF
C926 ffipg_3/ffi_0/q ffipg_3/ffi_0/qbar 0.32fF
C927 ffipg_3/ffi_0/inv_0/op gnd 0.27fF
C928 gnd ffipg_3/ffi_1/q 2.24fF
C929 ffipg_2/ffi_1/nand_3/a gnd 0.33fF
C930 gnd inv_5/w_0_6# 0.42fF
C931 gnd x4in 0.22fF
C932 gnd ffipg_0/ffi_0/inv_1/op 1.85fF
C933 sumffo_2/xor_0/w_n3_4# gnd 0.12fF
C934 sumffo_2/xor_0/inv_0/op gnd 0.32fF
C935 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_4/w_0_0# 0.06fF
C936 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/qbar 0.06fF
C937 y3in ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C938 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/q 0.31fF
C939 gnd ffo_0/d 0.45fF
C940 gnd sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C941 sumffo_0/ffo_0/inv_1/w_0_6# gnd 0.06fF
C942 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C943 ffipg_2/ffi_1/q ffipg_2/ffi_1/nand_6/a 0.31fF
C944 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C945 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a 0.13fF
C946 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C947 nor_0/b ffi_0/q 0.32fF
C948 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_3/b 0.33fF
C949 nor_3/b inv_5/w_0_6# 0.17fF
C950 cla_0/n inv_1/in 0.02fF
C951 inv_5/in cla_0/n 0.13fF
C952 ffipg_0/ffi_1/nand_0/w_0_0# gnd 0.10fF
C953 ffo_0/nand_3/a gnd 0.49fF
C954 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C955 ffi_0/nand_0/w_0_0# gnd 0.10fF
C956 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C957 sumffo_2/xor_0/inv_0/w_0_6# gnd 0.09fF
C958 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d 0.04fF
C959 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b 0.13fF
C960 clk ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C961 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_3/w_0_0# 0.04fF
C962 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C963 ffi_0/nand_3/a gnd 0.33fF
C964 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C965 sumffo_0/ffo_0/nand_1/a gnd 0.44fF
C966 gnd inv_8/in 0.43fF
C967 cla_0/l cla_1/l 0.08fF
C968 ffipg_2/ffi_0/inv_0/w_0_6# gnd 0.06fF
C969 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/k 0.45fF
C970 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C971 cla_1/inv_0/w_0_6# gnd 0.06fF
C972 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C973 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/nand_1/a 0.00fF
C974 gnd ffipg_1/ffi_1/qbar 0.67fF
C975 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/inv_0/op 0.06fF
C976 ffi_0/nand_3/b ffi_0/nand_1/a 0.00fF
C977 ffipg_2/ffi_1/inv_1/w_0_6# gnd 0.06fF
C978 ffipg_1/ffi_1/nand_2/w_0_0# ffipg_1/ffi_1/nand_3/a 0.04fF
C979 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C980 sumffo_0/ffo_0/nand_6/w_0_0# z1o 0.06fF
C981 ffi_0/nand_3/b ffi_0/nand_1/b 0.32fF
C982 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C983 cla_1/l gnd 0.40fF
C984 clk ffipg_3/ffi_1/inv_0/op 0.32fF
C985 ffipg_1/pggen_0/nand_0/w_0_0# cla_0/l 0.04fF
C986 sumffo_3/ffo_0/inv_1/w_0_6# sumffo_3/ffo_0/nand_0/b 0.03fF
C987 ffipg_0/ffi_0/q nor_0/a 0.03fF
C988 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/ffi_1/q 0.06fF
C989 ffipg_0/ffi_1/nand_1/a ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C990 ffipg_3/pggen_0/xor_0/inv_1/op gnd 0.35fF
C991 ffipg_1/pggen_0/nand_0/w_0_0# gnd 0.10fF
C992 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/ffi_0/q 0.12fF
C993 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C994 ffo_0/nand_1/b ffo_0/nand_3/b 0.32fF
C995 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C996 ffipg_0/ffi_0/nand_3/w_0_0# ffipg_0/ffi_0/nand_1/b 0.04fF
C997 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C998 sumffo_0/sbar z1o 0.32fF
C999 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C1000 cla_0/inv_0/in cla_1/p0 0.02fF
C1001 ffipg_0/ffi_1/inv_1/op gnd 1.85fF
C1002 gnd z2o 0.80fF
C1003 inv_5/in cla_2/l 0.05fF
C1004 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_3/b 0.33fF
C1005 nor_0/w_0_0# nor_0/a 0.06fF
C1006 inv_2/w_0_6# nor_1/b 0.03fF
C1007 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# 0.04fF
C1008 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C1009 ffipg_3/ffi_0/nand_6/a ffipg_3/ffi_0/nand_4/w_0_0# 0.04fF
C1010 ffipg_3/ffi_0/q ffipg_3/k 0.07fF
C1011 ffipg_1/ffi_1/inv_0/w_0_6# ffipg_1/ffi_1/inv_0/op 0.03fF
C1012 ffipg_0/ffi_1/nand_6/w_0_0# ffipg_0/ffi_1/qbar 0.04fF
C1013 cla_1/nor_1/w_0_0# cla_0/l 0.09fF
C1014 clk sumffo_1/ffo_0/nand_1/b 0.45fF
C1015 ffo_0/inv_1/w_0_6# gnd 0.06fF
C1016 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1017 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/b 0.32fF
C1018 cla_1/nor_1/w_0_0# gnd 0.31fF
C1019 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C1020 gnd ffipg_2/ffi_0/nand_7/w_0_0# 0.10fF
C1021 ffipg_2/ffi_0/nand_7/a ffipg_2/ffi_0/nand_1/b 0.13fF
C1022 ffipg_1/ffi_0/inv_1/w_0_6# gnd 0.06fF
C1023 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C1024 gnd sumffo_1/ffo_0/nand_3/a 0.48fF
C1025 nor_0/b sumffo_1/xor_0/a_38_n43# 0.01fF
C1026 clk y3in 0.68fF
C1027 ffipg_0/ffi_1/nand_3/b gnd 0.74fF
C1028 gnd sumffo_1/ffo_0/nand_7/w_0_0# 0.10fF
C1029 y4in clk 0.64fF
C1030 ffipg_3/ffi_0/nand_1/w_0_0# ffipg_3/ffi_0/nand_3/b 0.04fF
C1031 gnd ffipg_0/ffi_1/nand_7/a 0.37fF
C1032 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C1033 cla_0/n cla_2/l 0.32fF
C1034 ffipg_0/ffi_0/nand_1/b ffipg_0/ffi_0/inv_1/op 0.45fF
C1035 ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C1036 sumffo_0/ffo_0/nand_6/a z1o 0.31fF
C1037 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_6/a 0.31fF
C1038 gnd ffi_0/nand_1/a 0.44fF
C1039 gnd ffi_0/nand_1/b 0.57fF
C1040 gnd ffipg_2/ffi_0/qbar 0.67fF
C1041 gnd sumffo_3/ffo_0/inv_0/op 0.52fF
C1042 y2in ffipg_1/ffi_0/inv_0/op 0.04fF
C1043 ffipg_1/ffi_0/nand_3/a ffipg_1/ffi_0/nand_2/w_0_0# 0.04fF
C1044 inv_9/in ffo_0/d 0.04fF
C1045 gnd nor_4/w_0_0# 0.15fF
C1046 sumffo_1/ffo_0/nand_6/a z2o 0.31fF
C1047 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C1048 gnd ffi_0/q 0.80fF
C1049 x2in ffipg_1/ffi_1/inv_1/op 0.01fF
C1050 ffo_0/nand_2/w_0_0# gnd 0.10fF
C1051 sumffo_1/ffo_0/nand_5/w_0_0# gnd 0.10fF
C1052 y2in gnd 0.22fF
C1053 ffipg_0/ffi_0/inv_1/w_0_6# gnd 0.06fF
C1054 ffipg_0/ffi_0/nand_3/a ffipg_0/ffi_0/nand_3/b 0.31fF
C1055 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C1056 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_0/op 0.32fF
C1057 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C1058 y1in clk 0.68fF
C1059 ffipg_2/ffi_0/nand_5/w_0_0# gnd 0.10fF
C1060 couto ffo_0/qbar 0.32fF
C1061 gnd ffi_0/nand_2/w_0_0# 0.10fF
C1062 ffipg_2/ffi_1/nand_1/b ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1063 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/a 0.06fF
C1064 gnd ffipg_0/ffi_1/qbar 0.67fF
C1065 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.32fF
C1066 z1o gnd 0.80fF
C1067 cla_1/l inv_3/w_0_6# 0.06fF
C1068 sumffo_1/xor_0/inv_1/op nor_0/b 0.04fF
C1069 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/inv_1/op 0.33fF
C1070 ffipg_2/ffi_0/inv_1/w_0_6# ffipg_2/ffi_0/inv_1/op 0.04fF
C1071 ffipg_2/ffi_0/nand_3/w_0_0# gnd 0.11fF
C1072 sumffo_3/xor_0/a_10_10# ffipg_3/k 0.12fF
C1073 ffipg_1/ffi_0/nand_6/w_0_0# ffipg_1/ffi_0/q 0.06fF
C1074 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C1075 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C1076 gnd ffipg_2/ffi_1/nand_3/b 0.74fF
C1077 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_6/a 0.13fF
C1078 gnd ffipg_1/ffi_1/inv_0/op 0.27fF
C1079 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C1080 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C1081 cla_1/nor_1/w_0_0# cla_1/inv_0/in 0.05fF
C1082 clk ffipg_2/ffi_0/inv_0/op 0.32fF
C1083 ffipg_1/ffi_1/nand_1/b ffipg_1/ffi_1/inv_1/op 0.45fF
C1084 ffipg_1/ffi_1/nand_3/w_0_0# ffipg_1/ffi_1/nand_3/b 0.06fF
C1085 y4in ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1086 gnd ffipg_1/ffi_1/nand_3/a 0.33fF
C1087 cinin ffi_0/nand_2/w_0_0# 0.06fF
C1088 ffipg_2/ffi_1/nand_7/a gnd 0.37fF
C1089 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/qbar 0.00fF
C1090 ffipg_3/ffi_0/nand_0/w_0_0# clk 0.06fF
C1091 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_0/q 0.20fF
C1092 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C1093 sumffo_0/ffo_0/nand_7/w_0_0# z1o 0.04fF
C1094 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_1/w_0_6# 0.03fF
C1095 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/a 0.06fF
C1096 gnd ffipg_0/ffi_0/qbar 0.67fF
C1097 inv_7/w_0_6# inv_7/in 0.10fF
C1098 nand_2/b nor_0/b 0.04fF
C1099 ffipg_3/ffi_1/nand_2/w_0_0# x4in 0.06fF
C1100 nor_0/b ffi_0/nand_7/w_0_0# 0.06fF
C1101 clk ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C1102 inv_2/in nor_1/b 0.04fF
C1103 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op 0.06fF
C1104 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/qbar 0.31fF
C1105 ffipg_1/ffi_1/nand_2/w_0_0# x2in 0.06fF
C1106 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C1107 ffipg_0/ffi_0/q ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C1108 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/ffi_1/q 0.27fF
C1109 ffipg_3/ffi_0/nand_3/w_0_0# ffipg_3/ffi_0/nand_3/b 0.06fF
C1110 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C1111 gnd sumffo_1/ffo_0/nand_3/w_0_0# 0.11fF
C1112 ffipg_1/ffi_0/nand_6/a ffipg_1/ffi_0/qbar 0.00fF
C1113 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/w_0_0# 0.04fF
C1114 ffipg_3/ffi_0/q ffipg_3/pggen_0/xor_0/inv_0/op 0.20fF
C1115 clk ffo_0/nand_1/b 0.45fF
C1116 gnd sumffo_3/ffo_0/nand_7/a 0.33fF
C1117 sumffo_1/sbar z2o 0.32fF
C1118 ffipg_2/ffi_1/nand_1/a gnd 0.44fF
C1119 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/inv_0/w_0_6# 0.03fF
C1120 y4in ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C1121 inv_4/in gnd 0.33fF
C1122 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C1123 ffo_0/nand_0/b ffo_0/inv_0/op 0.32fF
C1124 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C1125 ffipg_2/ffi_1/inv_0/op ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C1126 sumffo_1/xor_0/inv_1/op ffipg_1/k 0.06fF
C1127 cla_2/nor_0/w_0_0# gnd 0.31fF
C1128 inv_8/w_0_6# nor_0/b 0.06fF
C1129 sumffo_2/xor_0/w_n3_4# inv_1/op 0.06fF
C1130 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C1131 ffipg_2/ffi_1/nand_1/a ffipg_2/ffi_1/nand_0/w_0_0# 0.04fF
C1132 inv_9/in nor_4/w_0_0# 0.11fF
C1133 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_6/a 0.31fF
C1134 gnd ffi_0/inv_0/op 0.27fF
C1135 ffipg_1/ffi_1/nand_5/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C1136 gnd ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C1137 ffo_0/nand_0/w_0_0# ffo_0/nand_1/a 0.04fF
C1138 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/sbar 0.06fF
C1139 nor_0/b inv_2/w_0_6# 0.06fF
C1140 cla_2/g1 cla_2/n 0.13fF
C1141 clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C1142 gnd ffipg_1/ffi_0/nand_2/w_0_0# 0.10fF
C1143 nor_1/w_0_0# gnd 0.15fF
C1144 ffipg_3/ffi_0/nand_6/w_0_0# gnd 0.10fF
C1145 x2in ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C1146 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1147 gnd ffipg_0/ffi_1/nand_3/w_0_0# 0.11fF
C1148 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C1149 nor_0/w_0_0# inv_0/op 0.10fF
C1150 ffipg_0/ffi_0/inv_0/op y1in 0.04fF
C1151 cla_2/inv_0/in cla_2/p1 0.02fF
C1152 ffipg_3/ffi_0/q ffipg_3/ffi_0/nand_6/a 0.31fF
C1153 clk ffipg_1/ffi_1/nand_1/a 0.13fF
C1154 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C1155 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C1156 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C1157 ffipg_1/pggen_0/nor_0/w_0_0# cla_1/p0 0.05fF
C1158 ffipg_0/ffi_1/inv_0/op clk 0.32fF
C1159 ffipg_0/ffi_0/nand_2/w_0_0# ffipg_0/ffi_0/nand_3/a 0.04fF
C1160 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C1161 sumffo_2/xor_0/inv_0/w_0_6# inv_1/op 0.06fF
C1162 ffi_0/nand_3/w_0_0# ffi_0/nand_3/a 0.06fF
C1163 sumffo_1/xor_0/inv_1/op gnd 0.35fF
C1164 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C1165 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b 0.13fF
C1166 inv_3/in gnd 0.47fF
C1167 ffipg_3/ffi_0/inv_1/op clk 0.07fF
C1168 ffipg_3/ffi_0/q ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C1169 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1170 ffipg_1/ffi_1/nand_7/w_0_0# ffipg_1/ffi_1/qbar 0.06fF
C1171 ffipg_1/k ffipg_1/ffi_0/q 0.07fF
C1172 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C1173 cla_0/l cla_2/p0 0.44fF
C1174 ffipg_3/ffi_0/nand_7/w_0_0# ffipg_3/ffi_0/q 0.04fF
C1175 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/inv_0/op 0.03fF
C1176 nand_2/b ffipg_1/k 0.15fF
C1177 cla_2/p0 gnd 1.06fF
C1178 ffo_0/nand_4/w_0_0# clk 0.06fF
C1179 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_0/op 0.32fF
C1180 nor_0/b sumffo_3/xor_0/w_n3_4# 0.01fF
C1181 cinin ffi_0/inv_0/op 0.04fF
C1182 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b 0.32fF
C1183 clk ffipg_0/ffi_0/nand_3/a 0.13fF
C1184 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_0/op 0.08fF
C1185 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C1186 ffipg_1/ffi_1/q ffipg_1/k 0.46fF
C1187 gnd ffipg_3/ffi_1/nand_6/a 0.37fF
C1188 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/q 0.00fF
C1189 inv_4/in cla_1/n 0.02fF
C1190 nor_0/a nor_0/b 0.32fF
C1191 ffo_0/nand_7/a gnd 0.33fF
C1192 gnd sumffo_3/ffo_0/nand_2/w_0_0# 0.10fF
C1193 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a 0.13fF
C1194 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C1195 cla_0/g0 nand_2/b 0.13fF
C1196 cla_0/l ffipg_1/ffi_0/q 0.13fF
C1197 clk ffo_0/nand_3/b 0.33fF
C1198 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/inv_1/op 0.06fF
C1199 ffi_0/nand_7/a ffi_0/nand_5/w_0_0# 0.04fF
C1200 cla_0/l nand_2/b 0.06fF
C1201 gnd ffipg_1/ffi_0/q 3.00fF
C1202 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b 0.32fF
C1203 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1204 cla_2/g1 cla_2/inv_0/op 0.35fF
C1205 cla_0/l ffipg_2/k 0.10fF
C1206 sumffo_2/xor_0/a_38_n43# nor_0/b 0.01fF
C1207 cla_2/g1 ffipg_3/ffi_0/q 0.13fF
C1208 ffipg_0/ffi_1/nand_0/w_0_0# ffipg_0/ffi_1/nand_1/a 0.04fF
C1209 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_0/inv_1/op 0.75fF
C1210 nand_2/b gnd 1.90fF
C1211 gnd ffipg_3/ffi_1/nand_0/w_0_0# 0.10fF
C1212 gnd ffi_0/nand_7/w_0_0# 0.10fF
C1213 gnd ffipg_0/ffi_0/nand_1/a 0.44fF
C1214 cla_2/p1 ffipg_3/ffi_1/q 0.22fF
C1215 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C1216 ffipg_2/ffi_1/nand_3/w_0_0# ffipg_2/ffi_1/nand_3/b 0.06fF
C1217 gnd ffipg_1/ffi_0/nand_1/a 0.44fF
C1218 gnd sumffo_3/ffo_0/nand_1/b 0.57fF
C1219 ffipg_2/k gnd 0.58fF
C1220 ffi_0/inv_1/op ffi_0/nand_3/b 0.33fF
C1221 ffipg_0/ffi_0/q ffipg_0/ffi_0/nand_7/a 0.00fF
C1222 ffipg_3/ffi_1/nand_4/w_0_0# ffipg_3/ffi_1/nand_6/a 0.04fF
C1223 ffipg_2/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1224 ffipg_1/ffi_1/q gnd 2.24fF
C1225 gnd sumffo_3/ffo_0/nand_0/b 0.53fF
C1226 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/k 0.02fF
C1227 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_3/b 0.31fF
C1228 ffipg_0/ffi_0/nand_4/w_0_0# gnd 0.10fF
C1229 cla_0/l ffipg_2/ffi_0/q 0.13fF
C1230 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1231 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C1232 x2in gnd 0.22fF
C1233 inv_8/w_0_6# gnd 0.15fF
C1234 gnd ffi_0/inv_0/w_0_6# 0.06fF
C1235 ffi_0/nand_3/w_0_0# ffi_0/nand_1/b 0.04fF
C1236 gnd ffipg_2/ffi_0/q 3.00fF
C1237 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C1238 cla_0/l inv_2/w_0_6# 0.06fF
C1239 nor_0/b sumffo_1/xor_0/a_10_10# 0.04fF
C1240 ffipg_0/ffi_0/nand_7/w_0_0# ffipg_0/ffi_0/qbar 0.06fF
C1241 cla_0/n cla_0/nand_0/w_0_0# 0.04fF
C1242 clk ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C1243 gnd inv_2/w_0_6# 0.17fF
C1244 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_0/nand_5/w_0_0# 0.06fF
C1245 ffipg_0/ffi_1/q ffipg_0/ffi_1/nand_7/a 0.00fF
C1246 ffipg_0/ffi_0/q ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1247 sumffo_0/ffo_0/nand_1/b clk 0.45fF
C1248 cla_1/inv_0/in cla_2/p0 0.02fF
C1249 inv_3/in inv_3/w_0_6# 0.10fF
C1250 inv_2/in nor_0/b 0.13fF
C1251 ffipg_2/ffi_1/inv_1/op ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C1252 ffipg_1/ffi_0/nand_1/b ffipg_1/ffi_0/nand_1/a 0.31fF
C1253 ffipg_0/ffi_0/nand_0/w_0_0# clk 0.06fF
C1254 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C1255 nor_0/a ffipg_1/k 0.06fF
C1256 ffipg_3/ffi_0/inv_1/op ffipg_3/ffi_1/inv_1/op 0.75fF
C1257 ffi_0/nand_6/a ffi_0/q 0.31fF
C1258 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_6/w_0_0# 0.04fF
C1259 ffipg_1/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C1260 nor_0/a ffipg_0/pggen_0/nor_0/w_0_0# 0.05fF
C1261 inv_4/in nor_2/b 0.16fF
C1262 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C1263 cla_0/l inv_7/in 0.13fF
C1264 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C1265 ffipg_3/ffi_1/inv_0/w_0_6# ffipg_3/ffi_1/inv_0/op 0.03fF
C1266 cinin ffi_0/inv_0/w_0_6# 0.06fF
C1267 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C1268 gnd inv_7/in 0.43fF
C1269 nor_0/a cla_0/g0 0.68fF
C1270 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/nand_1/a 0.00fF
C1271 nor_2/w_0_0# gnd 0.15fF
C1272 clk ffo_0/nand_6/a 0.13fF
C1273 clk sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C1274 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C1275 cla_1/nand_0/w_0_0# gnd 0.10fF
C1276 ffipg_1/ffi_1/nand_1/b gnd 0.57fF
C1277 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipg_1/ffi_0/q 0.23fF
C1278 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/ffi_1/q 0.06fF
C1279 ffi_0/inv_1/op gnd 1.89fF
C1280 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.35fF
C1281 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C1282 gnd sumffo_3/xor_0/w_n3_4# 0.12fF
C1283 ffipg_3/ffi_0/inv_1/w_0_6# ffipg_3/ffi_0/inv_1/op 0.04fF
C1284 ffi_0/nand_4/w_0_0# ffi_0/inv_1/op 0.06fF
C1285 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/k 0.01fF
C1286 nor_0/a cla_0/l 0.16fF
C1287 ffipg_0/ffi_1/q ffipg_0/ffi_1/qbar 0.32fF
C1288 ffipg_0/ffi_1/q ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C1289 nor_0/a gnd 0.54fF
C1290 ffipg_1/ffi_0/nand_7/a ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C1291 gnd nor_4/a 0.40fF
C1292 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_1/op 0.52fF
C1293 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/q 0.31fF
C1294 ffipg_0/ffi_1/inv_1/op ffipg_0/ffi_0/inv_1/op 0.75fF
C1295 ffipg_0/ffi_1/nand_6/w_0_0# ffipg_0/ffi_1/nand_6/a 0.06fF
C1296 inv_3/in nor_2/b 0.04fF
C1297 gnd ffo_0/nand_3/w_0_0# 0.11fF
C1298 sumffo_0/xor_0/inv_1/op nor_0/b 0.22fF
C1299 nand_2/b inv_3/w_0_6# 0.06fF
C1300 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/inv_1/op 0.06fF
C1301 ffipg_1/ffi_1/nand_1/w_0_0# gnd 0.10fF
C1302 ffipg_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C1303 ffipg_2/ffi_1/nand_5/w_0_0# gnd 0.10fF
C1304 gnd ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C1305 ffipg_0/ffi_1/nand_5/w_0_0# ffipg_0/ffi_1/nand_7/a 0.04fF
C1306 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/b 0.31fF
C1307 nor_0/a ffipg_0/k 0.05fF
C1308 ffi_0/inv_1/op ffi_0/inv_1/w_0_6# 0.04fF
C1309 nor_1/b inv_1/in 0.16fF
C1310 gnd sumffo_1/ffo_0/nand_2/a_13_n26# 0.01fF
C1311 sumffo_3/ffo_0/nand_6/a sumffo_3/sbar 0.00fF
C1312 gnd sumffo_3/sbar 0.62fF
C1313 cinin ffi_0/inv_1/op 0.01fF
C1314 cla_2/inv_0/w_0_6# gnd 0.06fF
C1315 cla_0/inv_0/op nand_2/b 0.09fF
C1316 ffipg_2/ffi_0/nand_1/a ffipg_2/ffi_0/nand_0/w_0_0# 0.04fF
C1317 clk sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C1318 clk ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C1319 ffipg_2/ffi_0/nand_4/w_0_0# gnd 0.10fF
C1320 gnd ffo_0/inv_0/op 0.37fF
C1321 ffipg_2/pggen_0/xor_0/inv_0/op gnd 0.32fF
C1322 ffipg_1/ffi_1/nand_5/w_0_0# gnd 0.10fF
C1323 sumffo_2/ffo_0/d clk 0.25fF
C1324 ffipg_3/ffi_1/nand_5/w_0_0# ffipg_3/ffi_1/nand_1/b 0.06fF
C1325 ffipg_2/ffi_1/nand_7/a ffipg_2/ffi_1/q 0.00fF
C1326 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k 0.52fF
C1327 cla_0/nor_1/w_0_0# cla_0/inv_0/in 0.05fF
C1328 nor_2/w_0_0# cla_1/n 0.06fF
C1329 cla_0/n nor_1/b 0.36fF
C1330 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C1331 ffipg_1/ffi_0/nand_1/w_0_0# ffipg_1/ffi_0/nand_1/a 0.06fF
C1332 gnd sumffo_1/xor_0/a_10_10# 0.93fF
C1333 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C1334 sumffo_0/ffo_0/nand_0/b gnd 0.58fF
C1335 gnd ffipg_2/ffi_0/inv_1/op 1.85fF
C1336 ffo_0/d nor_4/w_0_0# 0.03fF
C1337 y1in ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1338 gnd ffipg_0/ffi_0/nand_6/a 0.37fF
C1339 couto ffo_0/nand_7/a 0.00fF
C1340 sumffo_3/xor_0/a_10_10# sumffo_3/ffo_0/d 0.45fF
C1341 sumffo_1/ffo_0/nand_4/w_0_0# gnd 0.10fF
C1342 ffipg_0/ffi_0/inv_1/w_0_6# ffipg_0/ffi_0/inv_1/op 0.04fF
C1343 ffipg_2/k sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C1344 cla_1/inv_0/op cla_0/l 0.35fF
C1345 gnd ffipg_0/ffi_1/nand_6/a 0.37fF
C1346 ffo_0/nand_2/w_0_0# ffo_0/d 0.06fF
C1347 sumffo_2/ffo_0/nand_0/w_0_0# gnd 0.10fF
C1348 inv_2/in gnd 0.47fF
C1349 ffipg_3/ffi_1/nand_1/a ffipg_3/ffi_1/nand_0/w_0_0# 0.04fF
C1350 ffipg_2/ffi_0/nand_3/w_0_0# ffipg_2/ffi_0/nand_3/a 0.06fF
C1351 nor_1/w_0_0# inv_1/op 0.03fF
C1352 cla_1/inv_0/op gnd 0.27fF
C1353 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/nand_3/b 0.33fF
C1354 clk sumffo_3/ffo_0/d 0.04fF
C1355 ffi_0/nand_0/w_0_0# ffi_0/nand_1/a 0.04fF
C1356 ffipg_0/ffi_1/nand_3/a ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C1357 ffipg_0/ffi_0/inv_0/op ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C1358 ffipg_0/ffi_0/qbar ffipg_0/ffi_0/nand_6/w_0_0# 0.04fF
C1359 gnd ffipg_2/ffi_1/nand_6/w_0_0# 0.10fF
C1360 ffipg_1/pggen_0/xor_0/inv_1/op gnd 0.35fF
C1361 nor_0/a inv_0/in 0.02fF
C1362 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C1363 x1in ffipg_0/ffi_1/inv_0/op 0.04fF
C1364 clk ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1365 ffipg_2/ffi_1/nand_3/a ffipg_2/ffi_1/nand_3/b 0.31fF
C1366 ffipg_1/ffi_0/qbar ffipg_1/ffi_0/nand_7/a 0.31fF
C1367 sumffo_2/ffo_0/inv_0/op gnd 0.51fF
C1368 ffipg_1/ffi_1/nand_3/b ffipg_1/ffi_1/inv_1/op 0.33fF
C1369 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/inv_1/op 0.33fF
C1370 sumffo_2/sbar z3o 0.32fF
C1371 ffo_0/nand_5/w_0_0# ffo_0/nand_7/a 0.04fF
C1372 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_6/w_0_0# 0.04fF
C1373 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# 0.04fF
C1374 ffipg_2/ffi_0/nand_4/w_0_0# ffipg_2/ffi_0/nand_6/a 0.04fF
C1375 ffipg_1/ffi_0/qbar gnd 0.67fF
C1376 ffipg_0/ffi_1/nand_3/b ffipg_0/ffi_1/inv_1/op 0.33fF
C1377 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C1378 gnd ffipg_2/ffi_1/nand_4/w_0_0# 0.10fF
C1379 ffi_0/nand_3/a ffi_0/nand_2/w_0_0# 0.04fF
C1380 gnd ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C1381 gnd nor_3/w_0_0# 0.15fF
C1382 clk ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1383 inv_9/in nor_4/a 0.02fF
C1384 z4o sumffo_3/ffo_0/nand_7/a 0.00fF
C1385 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C1386 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C1387 sumffo_0/xor_0/inv_1/op gnd 0.35fF
C1388 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/nand_5/w_0_0# 0.04fF
C1389 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/inv_1/op 0.13fF
C1390 ffipg_1/ffi_1/nand_4/w_0_0# ffipg_1/ffi_1/nand_6/a 0.04fF
C1391 ffipg_0/ffi_0/nand_1/a ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1392 nor_2/w_0_0# nor_2/b 0.06fF
C1393 ffipg_2/ffi_0/nand_1/w_0_0# ffipg_2/ffi_0/nand_1/b 0.06fF
C1394 ffipg_1/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1395 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C1396 nor_3/b nor_3/w_0_0# 0.06fF
C1397 inv_6/in gnd 0.33fF
C1398 gnd ffipg_3/ffi_1/inv_0/op 0.27fF
C1399 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C1400 ffipg_3/ffi_1/inv_1/op ffipg_3/ffi_1/inv_1/w_0_6# 0.04fF
C1401 ffipg_1/ffi_1/nand_6/a ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C1402 clk ffipg_3/ffi_1/inv_1/op 0.07fF
C1403 ffipg_2/ffi_0/nand_7/w_0_0# ffipg_2/ffi_0/qbar 0.06fF
C1404 cla_2/p0 ffipg_2/ffi_1/q 0.22fF
C1405 ffipg_0/ffi_1/inv_0/op ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C1406 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C1407 ffipg_2/k inv_1/op 0.09fF
C1408 sumffo_0/xor_0/inv_0/op nor_0/b 0.20fF
C1409 cla_2/p1 cla_2/nor_0/w_0_0# 0.06fF
C1410 ffipg_2/ffi_0/nand_3/b ffipg_2/ffi_0/nand_1/b 0.32fF
C1411 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/ffi_0/q 0.23fF
C1412 ffipg_1/ffi_1/q ffipg_1/ffi_1/nand_7/w_0_0# 0.04fF
C1413 gnd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C1414 inv_6/in nor_3/b 0.16fF
C1415 sumffo_3/ffo_0/nand_3/w_0_0# gnd 0.11fF
C1416 sumffo_1/xor_0/inv_0/w_0_6# gnd 0.09fF
C1417 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C1418 inv_0/op cla_0/g0 0.34fF
C1419 ffipg_0/ffi_0/inv_0/op clk 0.32fF
C1420 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C1421 cla_0/g0 cla_0/inv_0/in 0.16fF
C1422 gnd ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C1423 gnd ffipg_3/ffi_0/qbar 0.67fF
C1424 ffi_0/nand_1/a ffi_0/nand_1/b 0.31fF
C1425 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C1426 sumffo_1/ffo_0/nand_1/b gnd 0.57fF
C1427 ffipg_3/ffi_0/inv_1/w_0_6# clk 0.06fF
C1428 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C1429 cla_0/l cla_0/inv_0/in 0.07fF
C1430 clk ffipg_1/ffi_0/inv_1/op 0.07fF
C1431 inv_0/op gnd 0.27fF
C1432 gnd y3in 0.22fF
C1433 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C1434 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1435 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/k 0.45fF
C1436 ffo_0/nand_0/b ffo_0/nand_1/a 0.13fF
C1437 cla_0/inv_0/in gnd 0.34fF
C1438 ffipg_2/k ffipg_2/ffi_1/q 0.46fF
C1439 ffipg_0/ffi_1/nand_7/a ffipg_0/ffi_1/qbar 0.31fF
C1440 y4in gnd 0.22fF
C1441 ffipg_0/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C1442 gnd ffipg_2/ffi_1/nand_7/w_0_0# 0.10fF
C1443 ffipg_2/ffi_1/nand_6/a ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C1444 sumffo_3/ffo_0/nand_4/w_0_0# clk 0.06fF
C1445 ffipg_1/ffi_0/nand_0/w_0_0# clk 0.06fF
C1446 cla_2/p1 cla_2/p0 0.24fF
C1447 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C1448 ffo_0/nand_7/a ffo_0/qbar 0.31fF
C1449 ffipg_3/ffi_0/q ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C1450 ffi_0/nand_0/w_0_0# ffi_0/inv_0/op 0.06fF
C1451 cla_2/l inv_7/w_0_6# 0.06fF
C1452 ffipg_3/ffi_1/qbar ffipg_3/ffi_1/nand_6/w_0_0# 0.04fF
C1453 ffipg_1/ffi_1/nand_0/w_0_0# ffipg_1/ffi_1/nand_1/a 0.04fF
C1454 ffo_0/inv_0/w_0_6# gnd 0.07fF
C1455 ffipg_2/ffi_1/qbar ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C1456 ffipg_2/ffi_1/q ffipg_2/ffi_0/q 0.73fF
C1457 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C1458 ffipg_3/ffi_0/nand_7/a ffipg_3/ffi_0/qbar 0.31fF
C1459 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C1460 gnd inv_4/op 0.58fF
C1461 ffipg_3/ffi_1/nand_6/a ffipg_3/ffi_1/q 0.31fF
C1462 ffipg_1/ffi_1/nand_4/w_0_0# gnd 0.10fF
C1463 ffipg_1/pggen_0/xor_0/a_10_10# gnd 0.93fF
C1464 y1in gnd 0.22fF
C1465 ffo_0/nand_0/b ffo_0/nand_0/w_0_0# 0.06fF
C1466 sumffo_3/xor_0/inv_0/w_0_6# inv_4/op 0.06fF
C1467 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_3/b 0.04fF
C1468 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C1469 sumffo_0/xor_0/w_n3_4# nor_0/b 0.06fF
C1470 nor_0/b sumffo_0/xor_0/a_10_10# 0.12fF
C1471 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C1472 ffipg_3/ffi_1/nand_1/b ffipg_3/ffi_1/nand_3/b 0.32fF
C1473 clk ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C1474 ffipg_3/ffi_1/nand_7/a ffipg_3/ffi_1/qbar 0.31fF
C1475 ffi_0/inv_1/op ffi_0/nand_6/a 0.13fF
C1476 ffipg_2/ffi_0/nand_6/a ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1477 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1478 gnd ffipg_1/ffi_1/nand_6/w_0_0# 0.10fF
C1479 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/k 0.02fF
C1480 clk sumffo_1/ffo_0/nand_3/b 0.33fF
C1481 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C1482 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_1/a 0.04fF
C1483 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C1484 cla_1/nor_0/w_0_0# cla_1/p0 0.06fF
C1485 ffipg_2/ffi_0/nand_7/a gnd 0.37fF
C1486 gnd sumffo_3/xor_0/inv_0/op 0.32fF
C1487 cla_0/l ffipg_3/k 0.10fF
C1488 inv_7/op inv_7/w_0_6# 0.03fF
C1489 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C1490 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/xor_0/inv_0/op 0.03fF
C1491 sumffo_1/ffo_0/d clk 0.04fF
C1492 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C1493 sumffo_3/ffo_0/inv_1/w_0_6# clk 0.06fF
C1494 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C1495 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C1496 gnd ffipg_3/ffi_0/nand_0/a_13_n26# 0.01fF
C1497 gnd ffipg_3/k 0.61fF
C1498 gnd ffipg_3/ffi_0/nand_4/w_0_0# 0.10fF
C1499 gnd ffipg_2/ffi_0/inv_0/op 0.27fF
C1500 ffipg_2/ffi_1/q ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1501 nor_0/a ffipg_0/ffi_1/q 0.22fF
C1502 inv_0/op inv_0/in 0.04fF
C1503 sumffo_0/xor_0/inv_0/op gnd 0.32fF
C1504 cla_1/l cla_2/p0 0.02fF
C1505 ffipg_0/ffi_0/nand_4/w_0_0# ffipg_0/ffi_0/inv_1/op 0.06fF
C1506 ffipg_3/ffi_0/nand_0/w_0_0# gnd 0.10fF
C1507 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# 0.04fF
C1508 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C1509 gnd ffipg_0/ffi_0/nand_7/a 0.37fF
C1510 ffipg_1/ffi_0/nand_3/b ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C1511 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# 0.04fF
C1512 x1in clk 0.68fF
C1513 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C1514 ffipg_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C1515 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C1516 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C1517 ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1518 ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1519 ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1520 ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1521 ffipg_3/ffi_1/qbar Gnd 0.42fF
C1522 ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1523 ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1524 ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1525 ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1526 ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1527 ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1528 ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1529 ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1530 x4in Gnd 0.51fF
C1531 ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1532 ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1533 ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1534 ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1535 ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1536 ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1537 ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1538 ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1539 ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1540 ffipg_3/ffi_0/qbar Gnd 0.42fF
C1541 ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1542 ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1543 ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1544 ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1545 ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1546 ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1547 ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1548 ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1549 y4in Gnd 0.51fF
C1550 ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1551 ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1552 ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1553 ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C1554 ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1555 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1556 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1557 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1558 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1559 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1560 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1561 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1562 ffipg_3/ffi_0/q Gnd 2.68fF
C1563 ffipg_3/ffi_1/q Gnd 2.93fF
C1564 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1565 ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1566 ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1567 ffi_0/nand_7/a Gnd 0.30fF
C1568 ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1569 ffi_0/nand_6/a Gnd 0.30fF
C1570 ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1571 ffi_0/inv_1/op Gnd 0.89fF
C1572 ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1573 ffi_0/nand_3/b Gnd 0.43fF
C1574 ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1575 ffi_0/nand_3/a Gnd 0.30fF
C1576 ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1577 clk Gnd 15.22fF
C1578 cinin Gnd 0.51fF
C1579 ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1580 ffi_0/inv_0/op Gnd 0.26fF
C1581 ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1582 ffi_0/nand_1/a Gnd 0.30fF
C1583 ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1584 ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1585 ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1586 ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C1587 ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1588 ffipg_2/ffi_1/qbar Gnd 0.42fF
C1589 ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C1590 ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1591 ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C1592 ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1593 ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C1594 ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1595 ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C1596 ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1597 x3in Gnd 0.51fF
C1598 ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1599 ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C1600 ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1601 ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C1602 ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1603 ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1604 ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1605 ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C1606 ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1607 ffipg_2/ffi_0/qbar Gnd 0.42fF
C1608 ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C1609 ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1610 ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C1611 ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1612 ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C1613 ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1614 ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C1615 ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1616 y3in Gnd 0.51fF
C1617 ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1618 ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C1619 ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1620 ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C1621 ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1622 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1623 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1624 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1625 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1626 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1627 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1628 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1629 ffipg_2/ffi_0/q Gnd 2.68fF
C1630 ffipg_2/ffi_1/q Gnd 2.93fF
C1631 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1632 ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1633 ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1634 ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C1635 ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1636 ffipg_1/ffi_1/qbar Gnd 0.42fF
C1637 ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C1638 ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1639 ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C1640 ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1641 ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C1642 ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1643 ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C1644 ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1645 x2in Gnd 0.51fF
C1646 ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1647 ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C1648 ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1649 ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C1650 ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1651 ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1652 ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1653 ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C1654 ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1655 ffipg_1/ffi_0/qbar Gnd 0.42fF
C1656 ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C1657 ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1658 ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C1659 ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1660 ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C1661 ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1662 ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C1663 ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1664 y2in Gnd 0.43fF
C1665 ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1666 ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C1667 ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1668 ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C1669 ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1670 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1671 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1672 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1673 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1674 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1675 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1676 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1677 ffipg_1/ffi_0/q Gnd 2.68fF
C1678 ffipg_1/ffi_1/q Gnd 2.93fF
C1679 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1680 inv_9/in Gnd 0.23fF
C1681 nor_4/w_0_0# Gnd 1.81fF
C1682 ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1683 ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1684 ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C1685 ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1686 ffipg_0/ffi_1/qbar Gnd 0.42fF
C1687 ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C1688 ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1689 ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C1690 ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1691 ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C1692 ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1693 ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C1694 ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1695 x1in Gnd 0.39fF
C1696 ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1697 ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C1698 ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1699 ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C1700 ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1701 ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1702 ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1703 ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C1704 ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1705 ffipg_0/ffi_0/qbar Gnd 0.42fF
C1706 ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C1707 ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1708 ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C1709 ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1710 ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C1711 ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1712 ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C1713 ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1714 y1in Gnd 0.51fF
C1715 ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1716 ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C1717 ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1718 ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C1719 ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C1720 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C1721 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C1722 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C1723 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C1724 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1725 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C1726 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1727 ffipg_0/ffi_0/q Gnd 2.68fF
C1728 ffipg_0/ffi_1/q Gnd 2.93fF
C1729 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C1730 nor_4/a Gnd 0.34fF
C1731 inv_8/in Gnd 0.22fF
C1732 inv_8/w_0_6# Gnd 1.40fF
C1733 inv_7/in Gnd 0.22fF
C1734 inv_7/w_0_6# Gnd 1.40fF
C1735 inv_5/in Gnd 0.22fF
C1736 inv_5/w_0_6# Gnd 1.40fF
C1737 nor_3/b Gnd 1.17fF
C1738 cla_2/n Gnd 0.36fF
C1739 nor_4/b Gnd 0.32fF
C1740 inv_6/in Gnd 0.23fF
C1741 nor_3/w_0_0# Gnd 1.81fF
C1742 cla_1/n Gnd 0.36fF
C1743 inv_4/in Gnd 0.23fF
C1744 nor_2/w_0_0# Gnd 1.81fF
C1745 nor_2/b Gnd 1.11fF
C1746 inv_3/in Gnd 0.22fF
C1747 inv_3/w_0_6# Gnd 1.40fF
C1748 nor_1/b Gnd 0.91fF
C1749 inv_2/in Gnd 0.22fF
C1750 inv_2/w_0_6# Gnd 1.40fF
C1751 inv_1/in Gnd 0.23fF
C1752 nor_1/w_0_0# Gnd 1.81fF
C1753 inv_0/in Gnd 0.23fF
C1754 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1755 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1756 ffo_0/nand_7/a Gnd 0.30fF
C1757 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1758 ffo_0/qbar Gnd 0.42fF
C1759 ffo_0/nand_6/a Gnd 0.30fF
C1760 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1761 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1762 ffo_0/nand_3/b Gnd 0.43fF
C1763 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1764 ffo_0/nand_3/a Gnd 0.30fF
C1765 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1766 ffo_0/nand_0/b Gnd 0.63fF
C1767 ffo_0/d Gnd 0.41fF
C1768 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1769 ffo_0/inv_0/op Gnd 0.26fF
C1770 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1771 ffo_0/nand_1/a Gnd 0.30fF
C1772 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1773 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1774 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1775 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1776 ffipg_3/k Gnd 1.88fF
C1777 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1778 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1779 inv_4/op Gnd 1.37fF
C1780 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1781 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1782 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1783 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1784 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1785 sumffo_3/sbar Gnd 0.43fF
C1786 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1787 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1788 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1789 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1790 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1791 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1792 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1793 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1794 sumffo_3/ffo_0/d Gnd 0.64fF
C1795 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1796 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1797 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1798 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1799 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1800 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1801 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1802 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1803 nand_2/b Gnd 1.99fF
C1804 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1805 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1806 ffipg_1/k Gnd 2.03fF
C1807 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1808 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1809 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1810 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1811 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1812 sumffo_1/sbar Gnd 0.43fF
C1813 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1814 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1815 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1816 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1817 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1818 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1819 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1820 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1821 sumffo_1/ffo_0/d Gnd 0.64fF
C1822 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1823 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1824 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1825 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1826 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1827 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1828 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1829 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1830 ffipg_2/k Gnd 1.93fF
C1831 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1832 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1833 inv_1/op Gnd 1.37fF
C1834 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1835 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1836 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1837 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1838 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1839 sumffo_2/sbar Gnd 0.43fF
C1840 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1841 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1842 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1843 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1844 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1845 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1846 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1847 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1848 sumffo_2/ffo_0/d Gnd 0.64fF
C1849 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1850 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1851 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1852 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1853 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1854 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1855 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1856 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1857 nor_0/b Gnd 2.77fF
C1858 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1859 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1860 ffipg_0/k Gnd 1.89fF
C1861 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1862 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1863 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1864 gnd Gnd 75.34fF
C1865 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1866 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1867 sumffo_0/sbar Gnd 0.43fF
C1868 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1869 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1870 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1871 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1872 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1873 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1874 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1875 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1876 sumffo_0/ffo_0/d Gnd 0.64fF
C1877 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1878 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1879 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1880 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1881 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1882 cla_2/p1 Gnd 1.09fF
C1883 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1884 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1885 cla_2/inv_0/in Gnd 0.27fF
C1886 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1887 cla_2/g1 Gnd 0.59fF
C1888 cla_2/inv_0/op Gnd 0.26fF
C1889 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1890 cla_1/nor_1/w_0_0# Gnd 1.23fF
C1891 cla_1/l Gnd 0.30fF
C1892 cla_1/nor_0/w_0_0# Gnd 1.23fF
C1893 cla_1/inv_0/in Gnd 0.27fF
C1894 cla_1/inv_0/w_0_6# Gnd 0.58fF
C1895 cla_1/inv_0/op Gnd 0.26fF
C1896 cla_1/nand_0/w_0_0# Gnd 0.82fF
C1897 inv_7/op Gnd 0.26fF
C1898 cla_0/nor_1/w_0_0# Gnd 1.23fF
C1899 cla_0/nor_0/w_0_0# Gnd 1.23fF
C1900 cla_0/inv_0/in Gnd 0.27fF
C1901 cla_0/inv_0/w_0_6# Gnd 0.58fF
C1902 cla_0/inv_0/op Gnd 0.26fF
C1903 cla_0/nand_0/w_0_0# Gnd 0.82fF
C1904 cla_2/l Gnd 0.75fF
C1905 inv_0/op Gnd 0.23fF
C1906 nor_0/w_0_0# Gnd 2.63fF
