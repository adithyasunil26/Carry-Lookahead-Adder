* SPICE3 file created from ffipgarrcla.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 vdd nand_1/b inv_1/in inv_1/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_1/in cla_0/l vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_1/in nand_1/b nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_2/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_0/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_2/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# nand_5/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd inv_7/op inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in nand_5/a vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in inv_7/op nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_0/g0 ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_0/g0 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1059 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1060 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1061 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1062 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1063 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1064 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 nor_0/a ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1069 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 gnd ffipgarr_0/ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1071 nor_0/a ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1073 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1074 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1076 ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1077 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1078 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 ffipgarr_0/ffipg_0/ffi_0/nand_1/a clk ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1081 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1082 ffipgarr_0/ffipg_0/ffi_0/nand_3/a y1in vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 ffipgarr_0/ffipg_0/ffi_0/nand_3/a clk ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1084 ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1086 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1088 ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1089 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1090 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1094 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1096 ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1097 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1098 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1101 vdd ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1102 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1107 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1108 ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1109 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1110 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1112 ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1113 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1114 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 ffipgarr_0/ffipg_0/ffi_1/nand_1/a clk ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1117 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1118 ffipgarr_0/ffipg_0/ffi_1/nand_3/a x1in vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 ffipgarr_0/ffipg_0/ffi_1/nand_3/a clk ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1122 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1124 ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1125 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1126 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1128 ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1129 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1130 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1133 vdd ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1134 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1136 ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1137 vdd ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1138 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1140 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1141 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1145 vdd ffipgarr_0/ffipg_1/ffi_0/q cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1146 cla_1/g0 ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1153 sumffo_1/k ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1154 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1155 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1156 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op sumffo_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 cla_1/p0 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1161 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 gnd ffipgarr_0/ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1163 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1165 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1166 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1168 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1169 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1170 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ffipgarr_0/ffipg_1/ffi_0/nand_1/a clk ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1172 ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1173 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1174 ffipgarr_0/ffipg_1/ffi_0/nand_3/a y2in vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 ffipgarr_0/ffipg_1/ffi_0/nand_3/a clk ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1176 ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1177 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1178 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1181 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1182 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1184 ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1185 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1186 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1188 ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1189 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1190 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1192 ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1193 vdd ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1194 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1201 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1202 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1204 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1205 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1206 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipgarr_0/ffipg_1/ffi_1/nand_1/a clk ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1208 ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1209 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1210 ffipgarr_0/ffipg_1/ffi_1/nand_3/a x2in vdd ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 ffipgarr_0/ffipg_1/ffi_1/nand_3/a clk ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1212 ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1213 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1214 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1216 ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1217 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1218 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1221 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1222 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1224 ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1225 vdd ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1226 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1228 ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1229 vdd ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1230 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1232 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1233 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1235 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1236 ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1237 vdd ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1238 cla_2/g0 ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 cla_2/g0 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1240 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1241 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1245 sumffo_2/k ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1246 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1247 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1248 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op sumffo_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1253 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 gnd ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1255 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1257 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1258 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1260 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1261 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1262 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 ffipgarr_0/ffipg_2/ffi_0/nand_1/a clk ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1264 ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1265 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1266 ffipgarr_0/ffipg_2/ffi_0/nand_3/a y3in vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 ffipgarr_0/ffipg_2/ffi_0/nand_3/a clk ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1268 ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1269 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1270 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1272 ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1273 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1274 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1276 ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1277 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1278 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1280 ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1281 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1282 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1284 ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1285 vdd ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1286 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1288 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1289 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1293 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1294 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1297 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1298 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 ffipgarr_0/ffipg_2/ffi_1/nand_1/a clk ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1301 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1302 ffipgarr_0/ffipg_2/ffi_1/nand_3/a x3in vdd ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 ffipgarr_0/ffipg_2/ffi_1/nand_3/a clk ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1304 ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1305 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1306 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1308 ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1309 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1310 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1313 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1314 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1316 ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1317 vdd ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1318 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1320 ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1321 vdd ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1322 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1325 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1326 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1327 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1328 ffipgarr_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1329 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1330 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/a vdd ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipgarr_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 vdd clk ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/inv_0/op vdd ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 ffipgarr_0/ffi_0/nand_1/a clk ffipgarr_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipgarr_0/ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1337 vdd clk ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1338 ffipgarr_0/ffi_0/nand_3/a cinin vdd ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 ffipgarr_0/ffi_0/nand_3/a clk ffipgarr_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 ffipgarr_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1341 vdd ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1342 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/a vdd ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1344 ffipgarr_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1345 vdd ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1346 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_3/b vdd ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1348 ffipgarr_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1349 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1350 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/inv_1/op vdd ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1352 ffipgarr_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 vdd nand_1/b nor_0/b ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 nor_0/b ffipgarr_0/ffi_0/nand_6/a vdd ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 nor_0/b nand_1/b ffipgarr_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipgarr_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 vdd nor_0/b nand_1/b ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 nand_1/b ffipgarr_0/ffi_0/nand_7/a vdd ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 nand_1/b nor_0/b ffipgarr_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipgarr_0/ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1361 ffipgarr_0/ffi_0/inv_0/op cinin vdd ffipgarr_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1362 ffipgarr_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1363 ffipgarr_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 vdd ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 cla_2/g1 ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1369 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1370 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1371 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1373 sumffo_3/k ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1374 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1375 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1376 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1381 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 gnd ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1383 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1385 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1386 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipgarr_0/ffipg_3/ffi_0/nand_1/a clk ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipgarr_0/ffipg_3/ffi_0/nand_3/a y4in vdd ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipgarr_0/ffipg_3/ffi_0/nand_3/a clk ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 vdd ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1417 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1418 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1419 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1421 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1422 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1425 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1426 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1427 ffipgarr_0/ffipg_3/ffi_1/nand_1/a clk ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1428 ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1429 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1430 ffipgarr_0/ffipg_3/ffi_1/nand_3/a x4in vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 ffipgarr_0/ffipg_3/ffi_1/nand_3/a clk ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1433 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1434 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1436 ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1437 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1438 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1440 ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1441 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1442 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1443 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1444 ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1445 vdd ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1446 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1448 ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1449 vdd ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1450 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1451 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1452 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1453 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1455 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1456 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1457 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1458 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1459 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1460 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1461 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1463 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1465 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1467 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1469 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1470 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a vdd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op vdd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1479 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1480 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 vdd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a vdd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 vdd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b vdd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 sumffo_0/ffo_0/nand_7/a clk vdd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 vdd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a vdd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 vdd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 z1o sumffo_0/ffo_0/nand_7/a vdd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1503 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1504 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1505 sumffo_0/ffo_0/nand_0/b clk vdd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 sumffo_0/xor_0/inv_0/op sumffo_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1507 sumffo_0/xor_0/inv_0/op sumffo_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1508 sumffo_0/xor_0/inv_1/op nand_1/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1509 sumffo_0/xor_0/inv_1/op nand_1/b vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 vdd nand_1/b sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1511 sumffo_0/ffo_0/d nand_1/b sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1512 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1513 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1514 sumffo_0/xor_0/a_10_n43# sumffo_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1515 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 sumffo_0/xor_0/a_10_10# sumffo_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1520 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a vdd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1522 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1523 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1524 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op vdd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1527 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1528 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1529 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1530 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1531 vdd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1532 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a vdd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1534 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1535 vdd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1536 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b vdd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1538 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 sumffo_2/ffo_0/nand_7/a clk vdd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 vdd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a vdd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 vdd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 z3o sumffo_2/ffo_0/nand_7/a vdd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1551 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1552 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1553 sumffo_2/ffo_0/nand_0/b clk vdd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 sumffo_2/xor_0/inv_0/op sumffo_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1555 sumffo_2/xor_0/inv_0/op sumffo_2/k vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1556 sumffo_2/xor_0/inv_1/op inv_2/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1557 sumffo_2/xor_0/inv_1/op inv_2/op vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 vdd inv_2/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1559 sumffo_2/ffo_0/d inv_2/op sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1560 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1561 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1562 sumffo_2/xor_0/a_10_n43# sumffo_2/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 sumffo_2/xor_0/a_10_10# sumffo_2/k vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a vdd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1571 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1572 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op vdd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1573 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 vdd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a vdd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 vdd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b vdd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 sumffo_1/ffo_0/nand_7/a clk vdd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 vdd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a vdd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 vdd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 z2o sumffo_1/ffo_0/nand_7/a vdd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1599 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1600 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1601 sumffo_1/ffo_0/nand_0/b clk vdd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 sumffo_1/xor_0/inv_0/op sumffo_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1603 sumffo_1/xor_0/inv_0/op sumffo_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1604 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1605 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1607 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1608 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1609 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1610 sumffo_1/xor_0/a_10_n43# sumffo_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1611 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 sumffo_1/xor_0/a_10_10# sumffo_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1614 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a vdd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op vdd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 vdd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a vdd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 vdd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b vdd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 sumffo_3/ffo_0/nand_7/a clk vdd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 vdd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a vdd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1643 vdd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1644 z4o sumffo_3/ffo_0/nand_7/a vdd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1645 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1647 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1648 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1649 sumffo_3/ffo_0/nand_0/b clk vdd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 sumffo_3/xor_0/inv_0/op sumffo_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 sumffo_3/xor_0/inv_0/op sumffo_3/k vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 sumffo_3/xor_0/inv_1/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 sumffo_3/xor_0/inv_1/op inv_4/op vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 vdd inv_4/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 sumffo_3/ffo_0/d inv_4/op sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 sumffo_3/xor_0/a_10_n43# sumffo_3/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 sumffo_3/xor_0/a_10_10# sumffo_3/k vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1663 vdd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1664 ffo_0/nand_3/b ffo_0/nand_1/a vdd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1665 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1666 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 vdd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffo_0/nand_1/a ffo_0/inv_0/op vdd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 vdd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffo_0/nand_3/a ffo_0/d vdd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 vdd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffo_0/nand_1/b ffo_0/nand_3/a vdd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 vdd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffo_0/nand_6/a ffo_0/nand_3/b vdd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 vdd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffo_0/nand_7/a clk vdd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 vdd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffo_0/qbar ffo_0/nand_6/a vdd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 vdd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 couto ffo_0/nand_7/a vdd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1695 ffo_0/inv_0/op ffo_0/d vdd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1696 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1697 ffo_0/nand_0/b clk vdd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 nor_1/b inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 nor_1/b inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 inv_2/op inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1703 inv_2/op inv_2/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1704 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1705 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1706 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1707 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1708 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1709 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 inv_2/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1711 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 gnd nor_1/b inv_2/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1713 inv_2/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1714 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1715 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1716 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1717 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1719 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 nor_4/a inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1721 nor_4/a inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1723 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1724 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1725 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1726 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1727 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1728 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1729 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1730 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1731 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1732 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1733 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 nor_4/b inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 nor_4/b inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffo_0/d inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 cla_1/nand_0/w_0_0# cla_0/n 0.01fF
C1 inv_0/op nor_0/w_0_0# 0.03fF
C2 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C3 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.00fF
C4 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.04fF
C5 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C6 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C7 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C8 vdd sumffo_1/ffo_0/nand_3/a 0.30fF
C9 sumffo_0/ffo_0/nand_3/a gnd 0.03fF
C10 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# vdd 0.10fF
C11 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.04fF
C12 ffipgarr_0/ffipg_2/ffi_1/qbar gnd 0.34fF
C13 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C14 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.31fF
C15 clk vdd 12.20fF
C16 cla_2/p0 vdd 0.43fF
C17 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.07fF
C18 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C19 ffipgarr_0/ffipg_1/ffi_0/q sumffo_1/k 0.07fF
C20 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.31fF
C21 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C22 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q 0.03fF
C23 cla_0/inv_0/op vdd 0.17fF
C24 clk sumffo_1/ffo_0/nand_1/b 0.45fF
C25 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C26 ffipgarr_0/ffipg_3/ffi_1/nand_1/b gnd 0.26fF
C27 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.04fF
C28 x3in vdd 0.04fF
C29 ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd 0.14fF
C30 clk sumffo_3/ffo_0/d 0.26fF
C31 ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd 0.03fF
C32 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.75fF
C33 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C34 cla_1/g0 cla_2/p0 0.32fF
C35 nand_2/b sumffo_2/k 0.03fF
C36 vdd sumffo_3/ffo_0/nand_3/b 0.39fF
C37 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# vdd 0.10fF
C38 sumffo_2/k inv_2/op 0.09fF
C39 vdd ffo_0/nand_1/w_0_0# 0.10fF
C40 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# vdd 0.11fF
C41 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.06fF
C42 cla_0/inv_0/op cla_1/g0 0.35fF
C43 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C44 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C45 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C46 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C47 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# vdd 0.10fF
C48 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C49 cla_0/g0 gnd 0.94fF
C50 ffipgarr_0/ffi_0/nand_6/a vdd 0.30fF
C51 ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd 0.30fF
C52 ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd 0.30fF
C53 cinin gnd 0.19fF
C54 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q 0.27fF
C55 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k 0.52fF
C56 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in 0.04fF
C57 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.08fF
C58 vdd sumffo_1/ffo_0/nand_1/a 0.30fF
C59 ffipgarr_0/ffipg_0/ffi_1/nand_1/b vdd 0.31fF
C60 nand_2/b cla_0/l 0.46fF
C61 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C62 cla_0/l inv_2/op 0.06fF
C63 gnd ffo_0/qbar 0.34fF
C64 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C65 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.04fF
C66 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C67 y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C68 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.04fF
C69 gnd inv_2/in 0.24fF
C70 vdd inv_4/op 0.25fF
C71 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_1/b 0.31fF
C72 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/inv_0/w_0_6# 0.03fF
C73 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C74 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C75 ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd 0.10fF
C76 vdd cla_0/n 0.68fF
C77 gnd sumffo_1/ffo_0/inv_0/op 0.10fF
C78 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C79 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.07fF
C80 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C81 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# 0.04fF
C82 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C83 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.31fF
C84 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C85 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.06fF
C86 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.06fF
C87 vdd nor_4/w_0_0# 0.15fF
C88 nor_1/w_0_0# inv_2/op 0.03fF
C89 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C90 sumffo_0/ffo_0/d vdd 0.04fF
C91 cla_1/inv_0/op vdd 0.17fF
C92 gnd inv_7/in 0.13fF
C93 vdd ffo_0/nand_7/a 0.30fF
C94 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.04fF
C95 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.45fF
C96 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op vdd 0.15fF
C97 y1in ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.01fF
C98 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.31fF
C99 cla_1/g0 cla_0/n 0.13fF
C100 cla_0/l cla_2/g0 0.08fF
C101 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# vdd 0.10fF
C102 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C103 vdd sumffo_3/ffo_0/nand_1/w_0_0# 0.10fF
C104 sumffo_2/ffo_0/nand_1/w_0_0# vdd 0.10fF
C105 ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd 0.17fF
C106 nand_2/b ffipgarr_0/ffipg_0/ffi_0/q 0.90fF
C107 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C108 sumffo_1/sbar sumffo_1/ffo_0/nand_7/a 0.31fF
C109 sumffo_1/ffo_0/nand_6/a z2o 0.31fF
C110 vdd sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C111 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# vdd 0.06fF
C112 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C113 ffo_0/nand_0/b ffo_0/inv_1/w_0_6# 0.03fF
C114 sumffo_0/ffo_0/nand_0/w_0_0# vdd 0.10fF
C115 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.06fF
C116 cla_1/nand_0/w_0_0# vdd 0.10fF
C117 vdd inv_8/w_0_6# 0.66fF
C118 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C119 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_0/b 0.40fF
C120 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.04fF
C121 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op gnd 0.20fF
C122 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C123 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q 0.22fF
C124 gnd sumffo_3/ffo_0/nand_3/a 0.03fF
C125 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/k 0.06fF
C126 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# sumffo_2/k 0.01fF
C127 nand_2/b cla_1/nor_0/w_0_0# 0.01fF
C128 inv_7/op inv_7/w_0_6# 0.03fF
C129 gnd sumffo_3/ffo_0/nand_1/b 0.26fF
C130 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.06fF
C131 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op sumffo_2/k 0.06fF
C132 nor_3/w_0_0# nor_3/b 0.06fF
C133 nor_0/a nor_0/b 0.39fF
C134 gnd ffo_0/d 0.26fF
C135 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# clk 0.06fF
C136 ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd 0.03fF
C137 clk sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C138 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_3/a 0.04fF
C139 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_3/b 0.04fF
C140 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C141 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C142 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.31fF
C143 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# vdd 0.06fF
C144 ffipgarr_0/ffi_0/nand_4/w_0_0# vdd 0.10fF
C145 ffipgarr_0/ffi_0/nand_2/w_0_0# ffipgarr_0/ffi_0/nand_3/a 0.04fF
C146 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.13fF
C147 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op sumffo_1/k 0.06fF
C148 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C149 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.04fF
C150 ffipgarr_0/ffi_0/nand_1/a gnd 0.14fF
C151 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_1/a 0.04fF
C152 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/ffo_0/nand_6/a 0.06fF
C153 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C154 vdd sumffo_2/ffo_0/nand_7/a 0.30fF
C155 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.31fF
C156 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C157 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.06fF
C158 gnd cla_1/n 0.08fF
C159 nor_3/w_0_0# inv_6/in 0.11fF
C160 nor_0/a inv_0/in 0.02fF
C161 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d 0.04fF
C162 vdd sumffo_1/ffo_0/nand_4/w_0_0# 0.10fF
C163 ffipgarr_0/ffipg_3/ffi_1/nand_3/a gnd 0.03fF
C164 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# vdd 0.10fF
C165 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.04fF
C166 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C167 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.06fF
C168 cla_1/l gnd 0.18fF
C169 cla_1/p0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C170 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.00fF
C171 cla_0/nor_0/a_13_6# nand_1/b 0.01fF
C172 sumffo_0/xor_0/a_10_10# vdd 0.93fF
C173 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# vdd 0.06fF
C174 x1in ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C175 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# vdd 0.10fF
C176 ffipgarr_0/ffipg_0/ffi_0/nand_1/b vdd 0.31fF
C177 cla_0/nor_0/w_0_0# vdd 0.32fF
C178 cla_2/l gnd 0.36fF
C179 clk sumffo_1/ffo_0/nand_6/a 0.13fF
C180 ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd 0.34fF
C181 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C182 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C183 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# sumffo_0/k 0.21fF
C184 gnd inv_4/in 0.24fF
C185 vdd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C186 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C187 sumffo_0/sbar z1o 0.32fF
C188 ffipgarr_0/ffipg_3/ffi_1/q sumffo_3/k 0.46fF
C189 cla_2/g1 vdd 0.35fF
C190 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.31fF
C191 nand_2/b nor_0/a 1.53fF
C192 vdd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C193 ffipgarr_0/ffipg_3/ffi_0/inv_1/op vdd 1.63fF
C194 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.31fF
C195 x1in ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.01fF
C196 vdd sumffo_1/ffo_0/nand_1/b 0.31fF
C197 ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd 0.34fF
C198 ffipgarr_0/ffipg_2/ffi_0/q vdd 0.38fF
C199 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in 0.04fF
C200 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.06fF
C201 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C202 y3in gnd 0.19fF
C203 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op sumffo_2/k 0.52fF
C204 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# vdd 0.10fF
C205 ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd 0.03fF
C206 cla_1/g0 vdd 0.49fF
C207 clk ffo_0/nand_4/w_0_0# 0.06fF
C208 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C209 vdd sumffo_3/ffo_0/d 0.04fF
C210 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C211 cla_2/p1 gnd 0.69fF
C212 ffipgarr_0/ffi_0/nand_7/w_0_0# vdd 0.10fF
C213 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C214 clk sumffo_3/ffo_0/nand_0/b 0.04fF
C215 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C216 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk 0.07fF
C217 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C218 ffipgarr_0/ffipg_0/ffi_0/qbar vdd 0.33fF
C219 ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd 0.39fF
C220 ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd 0.34fF
C221 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C222 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C223 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.32fF
C224 nor_0/b nand_1/b 2.65fF
C225 x3in ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.01fF
C226 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.06fF
C227 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.04fF
C228 vdd ffo_0/nand_3/a 0.30fF
C229 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q 0.27fF
C230 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C231 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# x4in 0.06fF
C232 ffipgarr_0/ffipg_2/ffi_0/inv_0/op ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.03fF
C233 sumffo_2/xor_0/inv_1/w_0_6# vdd 0.06fF
C234 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# vdd 0.10fF
C235 ffo_0/nand_6/a ffo_0/qbar 0.00fF
C236 sumffo_3/sbar z4o 0.32fF
C237 ffo_0/nand_3/w_0_0# ffo_0/nand_3/b 0.06fF
C238 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/sbar 0.04fF
C239 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C240 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.06fF
C241 sumffo_3/xor_0/inv_0/op sumffo_3/k 0.27fF
C242 sumffo_0/ffo_0/nand_3/w_0_0# vdd 0.11fF
C243 y4in gnd 0.19fF
C244 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# vdd 0.11fF
C245 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in 0.04fF
C246 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.31fF
C247 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.06fF
C248 cla_0/g0 cla_1/p0 0.33fF
C249 cla_0/l sumffo_2/ffo_0/nand_1/a 0.15fF
C250 ffo_0/nand_1/w_0_0# ffo_0/nand_1/a 0.06fF
C251 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/inv_0/op 0.06fF
C252 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/a 0.06fF
C253 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.13fF
C254 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.31fF
C255 inv_7/op nand_5/a 0.37fF
C256 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C257 ffipgarr_0/ffi_0/nand_1/b vdd 0.31fF
C258 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_1/b 0.04fF
C259 ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd 1.63fF
C260 nor_3/w_0_0# nor_4/a 0.03fF
C261 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C262 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.75fF
C263 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# clk 0.06fF
C264 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C265 cla_1/l inv_3/w_0_6# 0.06fF
C266 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.08fF
C267 ffipgarr_0/ffipg_0/ffi_1/nand_3/a clk 0.13fF
C268 cla_0/l nor_0/a 0.16fF
C269 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/qbar 0.00fF
C270 sumffo_0/ffo_0/nand_1/a gnd 0.03fF
C271 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.04fF
C272 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.06fF
C273 cla_2/p0 sumffo_3/k 0.09fF
C274 gnd sumffo_1/ffo_0/nand_7/a 0.03fF
C275 clk sumffo_0/ffo_0/nand_0/b 0.04fF
C276 x4in gnd 0.19fF
C277 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# clk 0.06fF
C278 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C279 nand_0/w_0_0# vdd 0.10fF
C280 vdd inv_1/in 0.30fF
C281 cla_2/n nor_3/b 0.37fF
C282 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.33fF
C283 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.04fF
C284 cla_1/p0 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C285 y1in clk 0.70fF
C286 inv_7/op inv_8/in 0.13fF
C287 nor_0/b sumffo_0/k 0.09fF
C288 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.31fF
C289 ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd 0.39fF
C290 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C291 cla_0/n nor_1/b 0.37fF
C292 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C293 nand_1/b sumffo_0/xor_0/inv_1/op 0.22fF
C294 clk ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C295 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# sumffo_3/k 0.21fF
C296 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C297 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.00fF
C298 ffipgarr_0/ffipg_2/ffi_1/q vdd 1.35fF
C299 ffipgarr_0/ffipg_1/ffi_1/inv_0/op clk 0.32fF
C300 ffipgarr_0/ffipg_1/ffi_1/q vdd 1.33fF
C301 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op sumffo_1/k 0.52fF
C302 ffipgarr_0/ffipg_0/ffi_0/q nor_0/a 0.14fF
C303 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C304 inv_6/in cla_2/n 0.02fF
C305 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C306 vdd sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C307 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.13fF
C308 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# vdd 0.06fF
C309 ffipgarr_0/ffipg_2/ffi_0/nand_1/a clk 0.13fF
C310 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_1/q 0.73fF
C311 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# vdd 0.10fF
C312 ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd 0.03fF
C313 cla_1/nor_1/a_13_6# gnd 0.01fF
C314 cla_1/g0 ffipgarr_0/ffipg_2/ffi_1/q 0.93fF
C315 x1in clk 0.70fF
C316 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.45fF
C317 vdd sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C318 vdd inv_7/w_0_6# 0.20fF
C319 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_0/b 0.06fF
C320 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b 0.13fF
C321 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.06fF
C322 x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C323 ffipgarr_0/ffipg_1/ffi_1/nand_3/a clk 0.13fF
C324 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# sumffo_1/k 0.01fF
C325 nand_2/b inv_3/in 0.13fF
C326 cla_2/l inv_5/in 0.03fF
C327 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C328 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C329 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C330 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_6/a 0.04fF
C331 sumffo_3/k cla_0/n 0.05fF
C332 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_1/op 0.06fF
C333 inv_4/op sumffo_3/k 0.09fF
C334 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_7/a 0.04fF
C335 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C336 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C337 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# vdd 0.10fF
C338 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.31fF
C339 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C340 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/b 0.32fF
C341 sumffo_0/ffo_0/nand_3/b gnd 0.35fF
C342 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# vdd 0.10fF
C343 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# cla_2/g1 0.04fF
C344 x2in ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.01fF
C345 cla_0/l nand_1/b 0.36fF
C346 clk sumffo_1/ffo_0/nand_3/b 0.33fF
C347 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_3/b 0.31fF
C348 nor_4/w_0_0# inv_9/in 0.11fF
C349 vdd sumffo_1/ffo_0/nand_6/a 0.30fF
C350 sumffo_0/ffo_0/nand_6/a gnd 0.03fF
C351 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C352 cla_2/inv_0/in cla_2/p1 0.02fF
C353 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C354 cinin ffipgarr_0/ffi_0/inv_1/op 0.01fF
C355 nor_0/b gnd 0.59fF
C356 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C357 nor_2/w_0_0# cla_1/n 0.06fF
C358 vdd sumffo_3/ffo_0/nand_3/w_0_0# 0.11fF
C359 cla_1/p0 cla_1/l 0.16fF
C360 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C361 vdd ffo_0/nand_2/w_0_0# 0.10fF
C362 sumffo_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C363 ffipgarr_0/ffipg_1/ffi_1/qbar vdd 0.33fF
C364 ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd 0.22fF
C365 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# vdd 0.10fF
C366 nand_5/a inv_8/w_0_6# 0.06fF
C367 cla_0/l sumffo_2/ffo_0/nand_3/a 0.15fF
C368 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C369 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_3/a 0.04fF
C370 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C371 ffipgarr_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C372 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.13fF
C373 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C374 vdd ffo_0/nand_4/w_0_0# 0.10fF
C375 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C376 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# vdd 0.11fF
C377 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# sumffo_2/k 0.21fF
C378 clk ffo_0/nand_3/b 0.33fF
C379 ffipgarr_0/ffi_0/nand_7/a vdd 0.30fF
C380 ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd 1.63fF
C381 ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd 0.39fF
C382 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C383 nor_2/w_0_0# inv_4/in 0.11fF
C384 gnd inv_0/in 0.24fF
C385 vdd sumffo_3/ffo_0/nand_0/b 0.15fF
C386 sumffo_2/ffo_0/d gnd 0.37fF
C387 ffipgarr_0/ffipg_0/ffi_0/q nand_1/b 0.02fF
C388 ffipgarr_0/ffipg_0/ffi_1/q nor_0/b 1.27fF
C389 ffo_0/nand_6/w_0_0# couto 0.06fF
C390 sumffo_2/xor_0/inv_0/op vdd 0.15fF
C391 ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd 0.34fF
C392 cla_1/nor_0/a_13_6# vdd 0.01fF
C393 vdd ffo_0/nand_1/a 0.30fF
C394 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.04fF
C395 vdd sumffo_1/k 0.26fF
C396 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C397 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.06fF
C398 cla_0/l inv_3/in 0.06fF
C399 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_0/b 0.40fF
C400 sumffo_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C401 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_3/b 0.00fF
C402 clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C403 ffipgarr_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffi_0/nand_7/a 0.06fF
C404 vdd ffo_0/nand_0/w_0_0# 0.10fF
C405 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d 0.04fF
C406 inv_8/w_0_6# inv_8/in 0.10fF
C407 ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd 0.34fF
C408 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C409 ffipgarr_0/ffipg_2/ffi_1/nand_1/b gnd 0.26fF
C410 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# vdd 0.10fF
C411 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.04fF
C412 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C413 nand_2/b gnd 1.54fF
C414 vdd nor_1/b 0.35fF
C415 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C416 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C417 gnd inv_2/op 0.26fF
C418 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/ffo_0/nand_7/a 0.06fF
C419 x3in ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C420 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# clk 0.06fF
C421 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# vdd 0.10fF
C422 nand_2/b cla_0/nor_1/w_0_0# 0.02fF
C423 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.06fF
C424 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.04fF
C425 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C426 sumffo_0/xor_0/inv_1/op gnd 0.20fF
C427 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.04fF
C428 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# vdd 0.10fF
C429 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# sumffo_2/k 0.45fF
C430 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# vdd 0.11fF
C431 inv_3/in nor_2/b 0.04fF
C432 vdd sumffo_1/xor_0/inv_1/op 0.15fF
C433 nor_3/b inv_5/w_0_6# 0.03fF
C434 ffipgarr_0/ffipg_1/ffi_1/nand_1/a clk 0.13fF
C435 ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd 0.30fF
C436 cla_2/g0 gnd 0.32fF
C437 nand_5/a vdd 0.02fF
C438 vdd inv_1/w_0_6# 0.15fF
C439 ffo_0/inv_0/op ffo_0/d 0.04fF
C440 ffipgarr_0/ffipg_2/ffi_1/nand_3/a clk 0.13fF
C441 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.45fF
C442 vdd inv_9/in 0.09fF
C443 sumffo_0/ffo_0/nand_0/b vdd 0.15fF
C444 vdd sumffo_3/k 0.31fF
C445 gnd sumffo_2/k 0.35fF
C446 ffipgarr_0/ffipg_0/ffi_1/nand_3/b gnd 0.35fF
C447 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C448 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.06fF
C449 ffipgarr_0/ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C450 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_7/a 0.13fF
C451 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.06fF
C452 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# vdd 0.10fF
C453 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C454 ffipgarr_0/ffipg_0/ffi_0/q sumffo_0/k 0.07fF
C455 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C456 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C457 y1in vdd 0.04fF
C458 inv_0/op vdd 0.17fF
C459 cla_0/g0 clk 0.10fF
C460 vdd z4o 0.28fF
C461 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C462 gnd sumffo_3/ffo_0/nand_6/a 0.03fF
C463 z3o gnd 0.52fF
C464 cla_2/inv_0/w_0_6# vdd 0.06fF
C465 gnd cla_2/n 0.22fF
C466 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# gnd 0.00fF
C467 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C468 nor_0/a nand_1/b 0.26fF
C469 cinin clk 0.70fF
C470 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# vdd 0.10fF
C471 ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd 0.17fF
C472 vdd inv_8/in 0.30fF
C473 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.31fF
C474 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# gnd 0.00fF
C475 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C476 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.13fF
C477 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.06fF
C478 ffipgarr_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C479 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar 0.32fF
C480 ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd 0.22fF
C481 cla_0/l gnd 0.88fF
C482 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/b 0.31fF
C483 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op vdd 0.15fF
C484 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/inv_1/w_0_6# 0.04fF
C485 ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd 0.30fF
C486 inv_7/op inv_7/in 0.04fF
C487 inv_6/in nor_3/b 0.16fF
C488 nor_0/b nor_0/w_0_0# 0.06fF
C489 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C490 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C491 ffipgarr_0/ffipg_1/ffi_0/inv_0/op clk 0.32fF
C492 x1in vdd 0.04fF
C493 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C494 gnd ffo_0/nand_0/b 0.43fF
C495 cla_1/nor_1/w_0_0# cla_2/g0 0.02fF
C496 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C497 sumffo_0/ffo_0/inv_0/op vdd 0.17fF
C498 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# vdd 0.10fF
C499 ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd 0.30fF
C500 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# vdd 0.93fF
C501 nand_2/b inv_3/w_0_6# 0.06fF
C502 sumffo_2/ffo_0/nand_2/w_0_0# cla_0/n 0.13fF
C503 inv_1/in nor_1/b 0.04fF
C504 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C505 vdd sumffo_1/ffo_0/nand_7/w_0_0# 0.10fF
C506 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C507 ffipgarr_0/ffipg_3/ffi_1/nand_7/a gnd 0.03fF
C508 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op gnd 0.17fF
C509 ffipgarr_0/ffipg_1/ffi_1/q sumffo_1/k 0.46fF
C510 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C511 gnd nor_2/b 0.10fF
C512 nor_0/w_0_0# inv_0/in 0.11fF
C513 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C514 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_1/op 0.52fF
C515 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/k 0.06fF
C516 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C517 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C518 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.04fF
C519 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# nand_1/b 0.02fF
C520 vdd sumffo_1/ffo_0/nand_3/b 0.39fF
C521 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# vdd 0.10fF
C522 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C523 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.00fF
C524 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op vdd 0.15fF
C525 ffipgarr_0/ffipg_0/ffi_0/q gnd 2.63fF
C526 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C527 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.06fF
C528 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_1/a 0.04fF
C529 z1o vdd 0.28fF
C530 ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 0.22fF
C531 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b 0.32fF
C532 sumffo_2/xor_0/w_n3_4# vdd 0.12fF
C533 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_7/a 0.04fF
C534 ffipgarr_0/ffipg_3/ffi_0/q gnd 2.62fF
C535 ffipgarr_0/ffi_0/inv_0/w_0_6# vdd 0.06fF
C536 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C537 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_2/ffi_0/q 0.23fF
C538 inv_1/w_0_6# inv_1/in 0.10fF
C539 nor_0/a sumffo_0/k 0.05fF
C540 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_6/a 0.04fF
C541 sumffo_2/xor_0/inv_1/op inv_2/op 0.22fF
C542 vdd sumffo_2/sbar 0.28fF
C543 ffipgarr_0/ffipg_2/ffi_0/qbar vdd 0.33fF
C544 ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd 0.22fF
C545 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# vdd 0.10fF
C546 ffipgarr_0/ffipg_0/ffi_0/nand_6/a gnd 0.03fF
C547 nor_4/a nor_4/b 0.35fF
C548 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C549 ffipgarr_0/ffipg_3/ffi_0/nand_1/b vdd 0.31fF
C550 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/ffi_0/nand_0/w_0_0# 0.06fF
C551 ffipgarr_0/ffipg_1/ffi_1/nand_1/b gnd 0.26fF
C552 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_1/q 0.73fF
C553 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.45fF
C554 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar 0.32fF
C555 nand_0/w_0_0# inv_0/op 0.06fF
C556 inv_2/in cla_0/n 0.02fF
C557 vdd ffo_0/nand_3/b 0.39fF
C558 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/b 0.31fF
C559 sumffo_2/ffo_0/nand_0/b gnd 0.38fF
C560 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.13fF
C561 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C562 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# clk 0.06fF
C563 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# sumffo_1/k 0.02fF
C564 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# vdd 0.10fF
C565 ffo_0/qbar ffo_0/nand_7/a 0.31fF
C566 ffipgarr_0/ffi_0/nand_1/a clk 0.13fF
C567 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b 0.32fF
C568 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C569 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/ffo_0/nand_6/a 0.06fF
C570 sumffo_0/sbar sumffo_0/ffo_0/nand_7/w_0_0# 0.06fF
C571 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C572 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.32fF
C573 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.06fF
C574 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.04fF
C575 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.04fF
C576 sumffo_0/ffo_0/nand_4/w_0_0# vdd 0.10fF
C577 ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd 0.03fF
C578 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# vdd 0.06fF
C579 cla_0/l inv_3/w_0_6# 0.17fF
C580 clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.13fF
C581 cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C582 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.06fF
C583 cla_1/l cla_2/p0 0.02fF
C584 gnd couto 0.52fF
C585 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C586 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.31fF
C587 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op gnd 0.20fF
C588 sumffo_2/k sumffo_2/xor_0/inv_1/op 0.06fF
C589 sumffo_0/ffo_0/nand_6/w_0_0# vdd 0.10fF
C590 ffipgarr_0/ffipg_3/ffi_0/qbar vdd 0.33fF
C591 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op 0.06fF
C592 sumffo_2/ffo_0/nand_1/a gnd 0.06fF
C593 cla_2/nor_1/w_0_0# cla_2/g1 0.02fF
C594 cla_2/nor_1/w_0_0# vdd 0.31fF
C595 cla_2/g0 cla_2/inv_0/in 0.16fF
C596 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.06fF
C597 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.04fF
C598 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# vdd 0.10fF
C599 y2in ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C600 cla_2/l cla_2/p0 0.16fF
C601 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.00fF
C602 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# sumffo_0/k 0.02fF
C603 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C604 sumffo_0/ffo_0/nand_6/a sumffo_0/sbar 0.00fF
C605 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.31fF
C606 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.13fF
C607 gnd nor_4/b 0.67fF
C608 clk sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C609 sumffo_0/ffo_0/nand_3/a vdd 0.30fF
C610 clk ffipgarr_0/ffi_0/inv_1/w_0_6# 0.06fF
C611 ffipgarr_0/ffipg_2/ffi_1/qbar vdd 0.33fF
C612 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# vdd 0.10fF
C613 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.06fF
C614 nand_2/b cla_1/p0 2.00fF
C615 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C616 y2in ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.01fF
C617 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.13fF
C618 nor_0/a gnd 0.29fF
C619 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.31fF
C620 ffo_0/nand_0/w_0_0# ffo_0/nand_1/a 0.04fF
C621 sumffo_2/ffo_0/nand_2/w_0_0# vdd 0.10fF
C622 ffipgarr_0/ffipg_3/ffi_1/nand_1/b vdd 0.31fF
C623 ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd 0.30fF
C624 inv_3/w_0_6# nor_2/b 0.03fF
C625 gnd inv_5/w_0_6# 0.01fF
C626 nand_2/b ffipgarr_0/ffipg_1/ffi_0/q 0.32fF
C627 inv_6/in nor_4/a 0.04fF
C628 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C629 nand_1/b sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C630 cla_2/p0 cla_2/p1 0.24fF
C631 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op gnd 0.20fF
C632 ffipgarr_0/ffi_0/inv_0/op gnd 0.10fF
C633 ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd 0.30fF
C634 y3in clk 0.70fF
C635 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.04fF
C636 ffipgarr_0/ffipg_0/ffi_0/nand_3/a clk 0.13fF
C637 nand_1/b sumffo_0/k 0.41fF
C638 vdd sumffo_1/ffo_0/nand_1/w_0_0# 0.10fF
C639 x4in ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.04fF
C640 ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd 0.10fF
C641 ffo_0/d nor_4/w_0_0# 0.03fF
C642 vdd sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C643 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/d 0.06fF
C644 ffipgarr_0/ffipg_0/ffi_1/q nor_0/a 0.22fF
C645 gnd ffo_0/inv_0/w_0_6# 0.01fF
C646 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C647 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C648 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C649 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# gnd 0.00fF
C650 ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd 0.34fF
C651 ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd 0.14fF
C652 cla_0/g0 vdd 0.50fF
C653 cla_0/n cla_1/n 0.09fF
C654 cla_1/p0 sumffo_2/k 2.09fF
C655 gnd nor_3/b 0.10fF
C656 sumffo_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C657 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.32fF
C658 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C659 cinin vdd 0.04fF
C660 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.00fF
C661 vdd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C662 ffipgarr_0/ffi_0/nand_2/w_0_0# vdd 0.10fF
C663 nand_2/b cla_0/nand_0/w_0_0# 0.01fF
C664 clk y4in 0.64fF
C665 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C666 cla_0/g0 cla_1/g0 0.18fF
C667 cla_2/l cla_0/n 0.31fF
C668 vdd ffo_0/qbar 0.28fF
C669 gnd sumffo_1/sbar 0.34fF
C670 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C671 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C672 inv_1/w_0_6# nor_1/b 0.03fF
C673 ffipgarr_0/ffipg_1/ffi_0/nand_1/b gnd 0.26fF
C674 inv_4/op inv_4/in 0.04fF
C675 vdd inv_2/in 0.09fF
C676 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_0/op 0.06fF
C677 sumffo_2/xor_0/a_10_10# inv_2/op 0.12fF
C678 ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd 0.17fF
C679 gnd inv_6/in 0.24fF
C680 vdd sumffo_1/ffo_0/inv_0/op 0.17fF
C681 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C682 gnd sumffo_3/ffo_0/nand_1/a 0.03fF
C683 ffipgarr_0/ffi_0/nand_3/b gnd 0.35fF
C684 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.06fF
C685 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.06fF
C686 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# clk 0.06fF
C687 cla_0/l cla_1/p0 0.02fF
C688 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# vdd 0.11fF
C689 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C690 vdd inv_7/in 0.34fF
C691 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.45fF
C692 sumffo_0/ffo_0/nand_7/a gnd 0.03fF
C693 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/xor_0/inv_0/op 0.03fF
C694 clk x4in 0.70fF
C695 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.06fF
C696 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C697 cla_0/inv_0/in gnd 0.35fF
C698 nand_1/b gnd 0.86fF
C699 vdd sumffo_3/ffo_0/nand_6/w_0_0# 0.10fF
C700 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C701 ffipgarr_0/ffipg_1/ffi_0/qbar gnd 0.34fF
C702 ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd 0.03fF
C703 ffipgarr_0/ffipg_0/ffi_1/qbar gnd 0.34fF
C704 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_0/q 0.12fF
C705 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C706 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C707 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in 0.04fF
C708 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.04fF
C709 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op vdd 0.15fF
C710 nor_2/w_0_0# nor_2/b 0.06fF
C711 clk ffo_0/nand_5/w_0_0# 0.06fF
C712 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/inv_0/w_0_6# 0.03fF
C713 vdd sumffo_3/ffo_0/nand_3/a 0.30fF
C714 sumffo_2/ffo_0/nand_3/a gnd 0.03fF
C715 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar 0.32fF
C716 ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd 0.03fF
C717 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# vdd 0.10fF
C718 ffipgarr_0/ffipg_0/ffi_0/nand_3/b gnd 0.35fF
C719 ffipgarr_0/ffipg_0/ffi_1/q nand_1/b 0.02fF
C720 ffo_0/nand_7/w_0_0# couto 0.04fF
C721 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C722 vdd sumffo_3/ffo_0/nand_1/b 0.31fF
C723 sumffo_2/ffo_0/nand_1/b gnd 0.38fF
C724 ffipgarr_0/ffipg_2/ffi_0/nand_1/b gnd 0.26fF
C725 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.00fF
C726 cla_1/inv_0/in cla_2/g0 0.04fF
C727 vdd ffo_0/d 0.19fF
C728 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C729 vdd sumffo_1/xor_0/a_10_10# 0.93fF
C730 ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd 0.03fF
C731 ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd 0.34fF
C732 cla_0/nand_0/w_0_0# cla_0/l 0.15fF
C733 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar 0.32fF
C734 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b 0.32fF
C735 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# vdd 0.06fF
C736 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.33fF
C737 nand_0/w_0_0# cla_0/g0 0.06fF
C738 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d 0.04fF
C739 nor_0/a nor_0/w_0_0# 0.06fF
C740 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_0/op 0.06fF
C741 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_6/a 0.04fF
C742 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# vdd 0.10fF
C743 ffipgarr_0/ffi_0/nand_1/a vdd 0.30fF
C744 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.04fF
C745 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C746 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C747 gnd inv_3/in 0.36fF
C748 ffo_0/nand_6/a couto 0.31fF
C749 nand_1/b sumffo_0/xor_0/w_n3_4# 0.06fF
C750 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C751 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C752 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C753 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k 0.06fF
C754 vdd cla_1/n 0.28fF
C755 cla_0/g0 ffipgarr_0/ffipg_1/ffi_1/q 0.84fF
C756 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C757 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.00fF
C758 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.00fF
C759 vdd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C760 ffipgarr_0/ffi_0/nand_0/w_0_0# gnd 0.00fF
C761 ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd 0.30fF
C762 cla_1/l vdd 0.27fF
C763 clk sumffo_0/ffo_0/nand_3/b 0.33fF
C764 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/b 0.31fF
C765 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.13fF
C766 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.04fF
C767 ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd 0.14fF
C768 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# gnd 0.00fF
C769 sumffo_0/k gnd 0.41fF
C770 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/b 0.32fF
C771 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C772 gnd sumffo_3/ffo_0/inv_0/op 0.32fF
C773 clk sumffo_0/ffo_0/nand_6/a 0.13fF
C774 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.13fF
C775 cla_2/l vdd 0.40fF
C776 gnd sumffo_3/ffo_0/inv_0/w_0_6# 0.01fF
C777 gnd nor_4/a 0.15fF
C778 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.04fF
C779 inv_5/w_0_6# inv_5/in 0.10fF
C780 vdd inv_4/in 0.09fF
C781 sumffo_2/ffo_0/nand_5/w_0_0# vdd 0.10fF
C782 ffipgarr_0/ffi_0/inv_1/w_0_6# vdd 0.06fF
C783 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# vdd 0.10fF
C784 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# vdd 0.10fF
C785 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# vdd 0.10fF
C786 sumffo_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C787 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.04fF
C788 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.31fF
C789 ffipgarr_0/ffi_0/nand_6/w_0_0# nand_1/b 0.06fF
C790 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk 0.07fF
C791 ffipgarr_0/ffipg_0/ffi_1/q sumffo_0/k 1.58fF
C792 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C793 cla_2/p1 cla_2/g1 0.00fF
C794 ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C795 cla_2/p1 vdd 0.31fF
C796 y3in vdd 0.04fF
C797 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C798 ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd 0.30fF
C799 nor_3/b inv_5/in 0.04fF
C800 ffo_0/nand_6/w_0_0# ffo_0/nand_6/a 0.06fF
C801 ffo_0/nand_5/w_0_0# ffo_0/nand_7/a 0.04fF
C802 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C803 gnd sumffo_3/ffo_0/nand_7/a 0.03fF
C804 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# gnd 0.00fF
C805 x2in gnd 0.19fF
C806 cla_1/p0 nor_0/a 0.24fF
C807 ffo_0/inv_0/op ffo_0/nand_0/b 0.32fF
C808 clk ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C809 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.04fF
C810 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.04fF
C811 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.31fF
C812 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# vdd 0.11fF
C813 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.04fF
C814 ffipgarr_0/ffi_0/nand_6/a nor_0/b 0.00fF
C815 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/b 0.31fF
C816 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_0/b 0.06fF
C817 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_3/b 0.00fF
C818 sumffo_0/xor_0/w_n3_4# sumffo_0/k 0.06fF
C819 inv_7/w_0_6# inv_7/in 0.10fF
C820 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C821 y4in ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C822 nand_2/b cla_2/p0 0.00fF
C823 clk inv_2/op 1.02fF
C824 sumffo_3/ffo_0/nand_6/a sumffo_3/sbar 0.00fF
C825 y4in vdd 0.04fF
C826 ffipgarr_0/ffi_0/nand_1/w_0_0# vdd 0.10fF
C827 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.00fF
C828 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.03fF
C829 y4in ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.01fF
C830 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.31fF
C831 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.06fF
C832 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# vdd 0.11fF
C833 gnd ffo_0/nand_1/b 0.26fF
C834 vdd sumffo_1/ffo_0/inv_0/w_0_6# 0.08fF
C835 inv_3/in inv_3/w_0_6# 0.10fF
C836 cla_0/l sumffo_2/ffo_0/nand_0/w_0_0# 0.17fF
C837 cla_0/nor_1/w_0_0# gnd 0.01fF
C838 cla_2/nand_0/w_0_0# gnd 0.01fF
C839 cla_0/g0 sumffo_1/k 0.07fF
C840 clk ffo_0/inv_1/w_0_6# 0.06fF
C841 sumffo_2/ffo_0/nand_7/w_0_0# z3o 0.04fF
C842 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C843 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# vdd 0.06fF
C844 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.06fF
C845 cla_2/p0 cla_2/g0 0.15fF
C846 ffipgarr_0/ffipg_0/ffi_1/q gnd 0.94fF
C847 sumffo_0/ffo_0/nand_1/a vdd 0.30fF
C848 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a 0.13fF
C849 x4in vdd 0.04fF
C850 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_0/q 0.73fF
C851 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.31fF
C852 cla_2/p0 sumffo_2/k 0.05fF
C853 vdd sumffo_1/ffo_0/nand_7/a 0.30fF
C854 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C855 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a 0.13fF
C856 sumffo_2/ffo_0/nand_6/a gnd 0.03fF
C857 ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd 0.03fF
C858 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.04fF
C859 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# clk 0.06fF
C860 cla_1/nor_1/w_0_0# gnd 0.01fF
C861 clk sumffo_3/ffo_0/nand_6/a 0.13fF
C862 cla_1/p0 nand_1/b 0.00fF
C863 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_0/q 0.23fF
C864 cla_0/inv_0/in cla_1/p0 0.02fF
C865 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_3/a 0.06fF
C866 nand_2/b cla_0/n 0.05fF
C867 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# y2in 0.06fF
C868 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# sumffo_1/k 0.21fF
C869 inv_2/op cla_0/n 0.70fF
C870 inv_2/in nor_1/b 0.16fF
C871 vdd ffo_0/nand_5/w_0_0# 0.10fF
C872 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C873 cla_0/nor_0/a_13_6# vdd 0.01fF
C874 vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C875 sumffo_3/ffo_0/nand_3/w_0_0# sumffo_3/ffo_0/nand_1/b 0.04fF
C876 sumffo_3/ffo_0/nand_0/w_0_0# vdd 0.10fF
C877 ffipgarr_0/ffipg_3/ffi_1/qbar gnd 0.34fF
C878 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.04fF
C879 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# clk 0.06fF
C880 cla_0/l clk 0.12fF
C881 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk 0.07fF
C882 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C883 vdd nor_3/w_0_0# 0.17fF
C884 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C885 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.04fF
C886 ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd 0.34fF
C887 cla_2/l inv_7/w_0_6# 0.06fF
C888 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar 0.32fF
C889 gnd sumffo_1/ffo_0/d 0.37fF
C890 ffipgarr_0/ffi_0/nand_3/a gnd 0.03fF
C891 clk ffo_0/nand_0/b 0.04fF
C892 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C893 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.06fF
C894 ffo_0/nand_2/w_0_0# ffo_0/d 0.06fF
C895 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a 0.13fF
C896 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/b 0.32fF
C897 sumffo_0/ffo_0/nand_7/w_0_0# vdd 0.10fF
C898 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.32fF
C899 inv_0/op cla_0/g0 0.32fF
C900 sumffo_3/xor_0/w_n3_4# inv_4/op 0.06fF
C901 gnd inv_3/w_0_6# 0.01fF
C902 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/nand_0/b 0.06fF
C903 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_0/qbar 0.04fF
C904 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C905 y3in ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C906 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.04fF
C907 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# sumffo_2/k 0.02fF
C908 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C909 sumffo_0/sbar sumffo_0/ffo_0/nand_7/a 0.31fF
C910 sumffo_0/ffo_0/nand_6/w_0_0# z1o 0.06fF
C911 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# vdd 0.10fF
C912 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.06fF
C913 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C914 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.06fF
C915 cla_1/inv_0/op cla_2/g0 0.35fF
C916 sumffo_0/ffo_0/nand_3/b vdd 0.39fF
C917 x4in ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.01fF
C918 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# vdd 0.10fF
C919 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/b 0.31fF
C920 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.06fF
C921 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.33fF
C922 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C923 sumffo_0/ffo_0/nand_6/a vdd 0.30fF
C924 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C925 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# vdd 0.06fF
C926 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C927 ffo_0/inv_0/op ffo_0/inv_0/w_0_6# 0.03fF
C928 sumffo_2/ffo_0/nand_3/w_0_0# vdd 0.11fF
C929 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/nand_1/a 0.04fF
C930 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b 0.32fF
C931 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C932 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C933 nor_0/b vdd 0.90fF
C934 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.33fF
C935 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C936 y2in gnd 0.19fF
C937 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# vdd 0.10fF
C938 ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd 0.03fF
C939 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# cla_2/p1 0.24fF
C940 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# sumffo_0/k 0.01fF
C941 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk 0.07fF
C942 cla_1/nand_0/w_0_0# cla_2/g0 0.06fF
C943 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C944 nand_1/b sumffo_0/xor_0/inv_0/op 0.20fF
C945 ffipgarr_0/ffipg_3/ffi_1/nand_1/a gnd 0.14fF
C946 ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd 1.63fF
C947 cla_0/l cla_0/n 0.83fF
C948 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/nand_3/a 0.04fF
C949 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_3/b 0.04fF
C950 nor_0/b ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C951 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_1/qbar 0.04fF
C952 cla_1/nor_0/w_0_0# cla_2/p0 0.06fF
C953 vdd inv_0/in 0.09fF
C954 inv_4/op sumffo_3/xor_0/a_10_10# 0.12fF
C955 sumffo_2/ffo_0/d vdd 0.04fF
C956 cla_2/inv_0/in gnd 0.35fF
C957 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# vdd 0.10fF
C958 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C959 clk sumffo_2/ffo_0/nand_0/b 0.04fF
C960 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# vdd 0.10fF
C961 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C962 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/inv_1/op 0.33fF
C963 gnd inv_5/in 0.17fF
C964 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C965 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.06fF
C966 nor_1/w_0_0# cla_0/n 0.06fF
C967 ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd 0.35fF
C968 gnd ffo_0/nand_6/a 0.03fF
C969 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C970 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.06fF
C971 clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.13fF
C972 ffo_0/d inv_9/in 0.04fF
C973 cinin ffipgarr_0/ffi_0/inv_0/w_0_6# 0.06fF
C974 cla_0/n nor_2/b 0.22fF
C975 vdd inv_2/op 0.34fF
C976 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.04fF
C977 ffipgarr_0/ffipg_2/ffi_1/nand_1/b vdd 0.31fF
C978 nand_2/b vdd 0.82fF
C979 cla_0/l cla_1/nand_0/w_0_0# 0.08fF
C980 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C981 sumffo_1/sbar z2o 0.32fF
C982 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# vdd 0.11fF
C983 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.04fF
C984 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C985 nand_2/b cla_1/g0 1.65fF
C986 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C987 nor_0/a clk 0.13fF
C988 cla_1/p0 gnd 0.74fF
C989 vdd ffo_0/inv_1/w_0_6# 0.06fF
C990 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C991 sumffo_0/xor_0/inv_1/op vdd 0.15fF
C992 vdd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C993 sumffo_2/ffo_0/nand_7/a z3o 0.00fF
C994 sumffo_0/xor_0/inv_0/op sumffo_0/k 0.27fF
C995 cla_2/g0 cla_2/g1 0.13fF
C996 cla_2/g0 vdd 0.45fF
C997 ffipgarr_0/ffi_0/inv_0/op clk 0.32fF
C998 ffipgarr_0/ffipg_1/ffi_0/q gnd 2.58fF
C999 ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd 0.03fF
C1000 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C1001 ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd 0.39fF
C1002 vdd sumffo_2/k 0.29fF
C1003 sumffo_3/xor_0/w_n3_4# sumffo_3/ffo_0/d 0.02fF
C1004 sumffo_2/xor_0/inv_1/w_0_6# inv_2/op 0.23fF
C1005 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# y3in 0.06fF
C1006 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C1007 cla_2/g0 ffipgarr_0/ffipg_2/ffi_0/q 0.13fF
C1008 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.06fF
C1009 ffipgarr_0/ffipg_0/ffi_1/inv_0/op clk 0.32fF
C1010 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.06fF
C1011 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C1012 sumffo_2/ffo_0/nand_3/b gnd 0.52fF
C1013 clk sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1014 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C1015 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.04fF
C1016 ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd 0.22fF
C1017 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C1018 cla_1/g0 cla_2/g0 0.13fF
C1019 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C1020 ffipgarr_0/ffipg_2/ffi_0/q sumffo_2/k 0.07fF
C1021 cla_1/g0 sumffo_2/k 0.56fF
C1022 vdd sumffo_3/ffo_0/nand_6/a 0.30fF
C1023 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/sbar 0.04fF
C1024 vdd z3o 0.28fF
C1025 cla_2/g1 cla_2/n 0.13fF
C1026 vdd cla_2/n 0.28fF
C1027 clk ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.32fF
C1028 cla_2/p1 sumffo_3/k 0.05fF
C1029 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# sumffo_3/k 0.01fF
C1030 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.04fF
C1031 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# 0.04fF
C1032 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# vdd 0.06fF
C1033 ffipgarr_0/ffipg_1/ffi_0/nand_1/a clk 0.13fF
C1034 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# vdd 0.10fF
C1035 ffipgarr_0/ffipg_0/ffi_0/nand_7/a gnd 0.03fF
C1036 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# clk 0.06fF
C1037 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C1038 sumffo_0/ffo_0/nand_5/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1039 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.06fF
C1040 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C1041 sumffo_2/ffo_0/nand_1/a cla_0/n 0.08fF
C1042 sumffo_1/xor_0/w_n3_4# sumffo_1/ffo_0/d 0.02fF
C1043 sumffo_0/sbar gnd 0.34fF
C1044 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C1045 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# vdd 0.10fF
C1046 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.33fF
C1047 cla_0/nand_0/w_0_0# gnd 0.01fF
C1048 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_1/w_0_6# 0.03fF
C1049 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a 0.13fF
C1050 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# vdd 0.06fF
C1051 ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd 1.63fF
C1052 cla_0/l vdd 1.74fF
C1053 ffo_0/nand_7/a couto 0.00fF
C1054 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.06fF
C1055 vdd sumffo_3/xor_0/a_10_10# 0.93fF
C1056 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# vdd 0.93fF
C1057 vdd ffo_0/nand_0/b 0.15fF
C1058 gnd sumffo_1/ffo_0/nand_0/b 0.45fF
C1059 ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd 0.35fF
C1060 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C1061 clk sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C1062 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.06fF
C1063 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.06fF
C1064 nand_2/b inv_1/in 0.04fF
C1065 vdd nor_1/w_0_0# 0.15fF
C1066 vdd sumffo_1/xor_0/inv_0/op 0.15fF
C1067 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/a 0.06fF
C1068 sumffo_0/xor_0/inv_0/op gnd 0.17fF
C1069 ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd 0.03fF
C1070 nand_0/w_0_0# nand_2/b 0.04fF
C1071 nor_4/b nor_4/w_0_0# 0.06fF
C1072 sumffo_3/ffo_0/d sumffo_3/xor_0/a_10_10# 0.45fF
C1073 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C1074 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C1075 ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd 0.34fF
C1076 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op vdd 0.15fF
C1077 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.04fF
C1078 cla_0/inv_0/w_0_6# vdd 0.06fF
C1079 cla_0/n inv_5/w_0_6# 0.06fF
C1080 clk nand_1/b 0.05fF
C1081 clk sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C1082 vdd nor_2/b 0.35fF
C1083 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C1084 sumffo_2/ffo_0/nand_6/w_0_0# vdd 0.10fF
C1085 cla_2/nor_0/w_0_0# vdd 0.31fF
C1086 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# vdd 0.10fF
C1087 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.13fF
C1088 nand_2/b ffipgarr_0/ffipg_2/ffi_1/q 0.69fF
C1089 cinin ffipgarr_0/ffi_0/nand_2/w_0_0# 0.06fF
C1090 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.06fF
C1091 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_0/q 0.20fF
C1092 ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd 0.22fF
C1093 ffipgarr_0/ffipg_0/ffi_0/q vdd 0.38fF
C1094 cla_1/inv_0/in gnd 0.35fF
C1095 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C1096 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_3/b 0.00fF
C1097 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.06fF
C1098 ffipgarr_0/ffi_0/nand_3/w_0_0# vdd 0.11fF
C1099 ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.31fF
C1100 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/qbar 0.04fF
C1101 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C1102 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C1103 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1104 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# y4in 0.06fF
C1105 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1106 inv_8/w_0_6# nor_4/b 0.03fF
C1107 ffo_0/nand_0/b ffo_0/nand_3/a 0.13fF
C1108 ffipgarr_0/ffipg_3/ffi_0/q vdd 0.38fF
C1109 ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 0.13fF
C1110 ffipgarr_0/ffi_0/inv_1/op gnd 0.22fF
C1111 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# vdd 0.11fF
C1112 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.32fF
C1113 gnd ffo_0/inv_0/op 0.34fF
C1114 ffipgarr_0/ffipg_2/ffi_0/nand_3/a clk 0.13fF
C1115 ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd 0.15fF
C1116 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C1117 ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd 1.63fF
C1118 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/qbar 0.04fF
C1119 ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd 0.34fF
C1120 clk sumffo_2/ffo_0/nand_1/b 0.45fF
C1121 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.00fF
C1122 ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd 0.10fF
C1123 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# vdd 0.10fF
C1124 ffipgarr_0/ffipg_1/ffi_1/nand_1/b vdd 0.31fF
C1125 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar 0.32fF
C1126 cla_1/nor_0/w_0_0# vdd 0.32fF
C1127 vdd sumffo_1/ffo_0/nand_2/w_0_0# 0.10fF
C1128 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1129 nor_0/b ffipgarr_0/ffi_0/nand_7/a 0.31fF
C1130 ffipgarr_0/ffi_0/nand_6/a nand_1/b 0.31fF
C1131 sumffo_2/ffo_0/nand_0/b vdd 0.15fF
C1132 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C1133 ffipgarr_0/ffipg_3/ffi_1/q gnd 0.93fF
C1134 ffipgarr_0/ffipg_2/ffi_1/q sumffo_2/k 2.17fF
C1135 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/k 0.06fF
C1136 sumffo_3/sbar sumffo_3/ffo_0/nand_7/a 0.31fF
C1137 cla_2/inv_0/op gnd 0.10fF
C1138 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/qbar 0.00fF
C1139 ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd 0.30fF
C1140 sumffo_2/ffo_0/nand_4/w_0_0# cla_0/n 0.24fF
C1141 cla_0/l inv_1/in 0.08fF
C1142 vdd couto 0.28fF
C1143 gnd z2o 0.52fF
C1144 sumffo_1/ffo_0/d sumffo_1/ffo_0/nand_0/b 0.40fF
C1145 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.04fF
C1146 ffipgarr_0/ffi_0/nand_0/w_0_0# clk 0.06fF
C1147 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C1148 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op vdd 0.15fF
C1149 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op gnd 0.17fF
C1150 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C1151 clk ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1152 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C1153 ffipgarr_0/ffipg_0/ffi_0/nand_1/a clk 0.13fF
C1154 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op 0.06fF
C1155 sumffo_2/ffo_0/inv_0/op gnd 0.10fF
C1156 sumffo_2/ffo_0/nand_1/a vdd 0.30fF
C1157 ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd 0.10fF
C1158 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# 0.04fF
C1159 gnd sumffo_3/sbar 0.34fF
C1160 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C1161 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C1162 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C1163 ffipgarr_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.04fF
C1164 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C1165 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C1166 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# clk 0.06fF
C1167 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C1168 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# vdd 0.10fF
C1169 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.06fF
C1170 vdd nor_4/b 0.41fF
C1171 sumffo_2/ffo_0/nand_3/a cla_0/n 0.07fF
C1172 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C1173 clk ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C1174 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.45fF
C1175 ffipgarr_0/ffipg_0/ffi_0/inv_0/op gnd 0.10fF
C1176 nor_0/a vdd 0.29fF
C1177 sumffo_2/ffo_0/nand_1/b cla_0/n 0.05fF
C1178 sumffo_2/xor_0/inv_0/op inv_2/op 0.20fF
C1179 nand_2/b cla_1/nor_0/a_13_6# 0.01fF
C1180 inv_4/op sumffo_3/xor_0/inv_1/op 0.22fF
C1181 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C1182 nand_2/b sumffo_1/k 0.51fF
C1183 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op vdd 0.15fF
C1184 ffipgarr_0/ffi_0/inv_0/op vdd 0.17fF
C1185 ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd 0.03fF
C1186 cla_0/l inv_7/w_0_6# 0.06fF
C1187 vdd inv_5/w_0_6# 0.15fF
C1188 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.00fF
C1189 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# clk 0.06fF
C1190 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q 0.27fF
C1191 x2in clk 0.70fF
C1192 sumffo_0/ffo_0/nand_1/b gnd 0.26fF
C1193 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C1194 ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd 0.17fF
C1195 sumffo_0/ffo_0/nand_1/w_0_0# vdd 0.10fF
C1196 cla_0/n inv_3/in 0.02fF
C1197 vdd ffo_0/nand_6/w_0_0# 0.10fF
C1198 sumffo_0/ffo_0/inv_1/w_0_6# vdd 0.06fF
C1199 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar 0.32fF
C1200 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.04fF
C1201 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.06fF
C1202 cla_2/nor_1/a_13_6# gnd 0.01fF
C1203 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C1204 ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd 0.35fF
C1205 inv_7/op gnd 0.16fF
C1206 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q 0.21fF
C1207 vdd ffo_0/inv_0/w_0_6# 0.06fF
C1208 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C1209 ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd 0.17fF
C1210 ffipgarr_0/ffipg_1/ffi_1/inv_0/op ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.03fF
C1211 ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd 0.30fF
C1212 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# vdd 0.10fF
C1213 vdd nor_3/b 0.35fF
C1214 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.04fF
C1215 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# clk 0.06fF
C1216 clk gnd 8.12fF
C1217 cla_2/p0 gnd 0.74fF
C1218 gnd sumffo_1/ffo_0/nand_3/a 0.03fF
C1219 sumffo_2/xor_0/inv_0/op sumffo_2/k 0.27fF
C1220 inv_0/op inv_0/in 0.04fF
C1221 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C1222 vdd sumffo_1/sbar 0.28fF
C1223 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C1224 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.32fF
C1225 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C1226 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C1227 nand_2/b inv_1/w_0_6# 0.01fF
C1228 clk ffo_0/nand_1/b 0.45fF
C1229 x3in gnd 0.19fF
C1230 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# 0.04fF
C1231 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.04fF
C1232 ffipgarr_0/ffipg_1/ffi_0/nand_1/b vdd 0.31fF
C1233 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.16fF
C1234 cla_0/inv_0/op gnd 0.15fF
C1235 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.06fF
C1236 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.06fF
C1237 vdd inv_6/in 0.09fF
C1238 gnd sumffo_3/ffo_0/nand_3/b 0.35fF
C1239 sumffo_0/ffo_0/nand_7/w_0_0# z1o 0.04fF
C1240 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# vdd 0.11fF
C1241 cla_2/l inv_7/in 0.13fF
C1242 nand_1/b sumffo_0/xor_0/a_10_10# 0.12fF
C1243 sumffo_0/ffo_0/nand_5/w_0_0# vdd 0.10fF
C1244 ffipgarr_0/ffi_0/nand_3/b vdd 0.39fF
C1245 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C1246 nor_4/a nor_4/w_0_0# 0.06fF
C1247 vdd sumffo_3/ffo_0/nand_1/a 0.30fF
C1248 cla_0/nor_0/w_0_0# nand_1/b 0.01fF
C1249 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C1250 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.06fF
C1251 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.33fF
C1252 sumffo_0/ffo_0/nand_7/a vdd 0.30fF
C1253 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C1254 sumffo_2/ffo_0/nand_4/w_0_0# vdd 0.10fF
C1255 nand_1/b vdd 1.12fF
C1256 ffipgarr_0/ffi_0/nand_6/a gnd 0.03fF
C1257 ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd 0.14fF
C1258 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.13fF
C1259 ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd 0.03fF
C1260 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1261 cla_0/inv_0/in vdd 0.05fF
C1262 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C1263 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1264 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C1265 sumffo_3/xor_0/w_n3_4# sumffo_3/k 0.06fF
C1266 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C1267 sumffo_0/ffo_0/nand_6/a z1o 0.31fF
C1268 ffipgarr_0/ffipg_1/ffi_0/qbar vdd 0.33fF
C1269 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# vdd 0.10fF
C1270 cla_2/g0 sumffo_3/k 0.10fF
C1271 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C1272 ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd 0.34fF
C1273 ffipgarr_0/ffipg_0/ffi_1/qbar vdd 0.33fF
C1274 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.31fF
C1275 ffipgarr_0/ffipg_0/ffi_1/nand_1/b gnd 0.26fF
C1276 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.04fF
C1277 gnd sumffo_1/ffo_0/nand_1/a 0.27fF
C1278 cla_0/l nor_1/b 0.10fF
C1279 ffo_0/nand_1/a ffo_0/nand_0/b 0.13fF
C1280 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C1281 ffipgarr_0/ffi_0/nand_7/w_0_0# nand_1/b 0.04fF
C1282 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# clk 0.06fF
C1283 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# sumffo_1/k 0.45fF
C1284 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.32fF
C1285 cla_1/nor_1/w_0_0# cla_2/p0 0.06fF
C1286 cla_1/g0 cla_0/inv_0/in 0.04fF
C1287 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# vdd 0.10fF
C1288 sumffo_2/ffo_0/nand_0/a_13_n26# gnd 0.00fF
C1289 ffo_0/nand_0/w_0_0# ffo_0/nand_0/b 0.06fF
C1290 gnd inv_4/op 0.21fF
C1291 sumffo_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C1292 clk sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1293 sumffo_2/ffo_0/nand_3/a vdd 0.30fF
C1294 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C1295 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C1296 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C1297 ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd 0.30fF
C1298 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# clk 0.06fF
C1299 ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd 0.39fF
C1300 gnd cla_0/n 0.52fF
C1301 sumffo_2/ffo_0/nand_1/a_13_n26# gnd 0.01fF
C1302 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C1303 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1304 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.06fF
C1305 sumffo_2/ffo_0/nand_1/b vdd 0.31fF
C1306 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1307 ffipgarr_0/ffipg_2/ffi_0/nand_1/b vdd 0.31fF
C1308 clk sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C1309 sumffo_0/ffo_0/d gnd 0.37fF
C1310 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C1311 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# vdd 0.10fF
C1312 ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd 0.34fF
C1313 cla_1/inv_0/op gnd 0.15fF
C1314 nor_1/w_0_0# nor_1/b 0.06fF
C1315 vdd sumffo_3/xor_0/inv_1/op 0.15fF
C1316 clk sumffo_1/ffo_0/d 0.05fF
C1317 gnd ffo_0/nand_7/a 0.03fF
C1318 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1319 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C1320 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C1321 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C1322 ffipgarr_0/ffi_0/nand_3/a clk 0.13fF
C1323 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op gnd 0.20fF
C1324 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/qbar 0.00fF
C1325 cla_0/l inv_1/w_0_6# 0.28fF
C1326 sumffo_2/ffo_0/nand_1/w_0_0# gnd 0.00fF
C1327 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C1328 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C1329 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.75fF
C1330 ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd 0.10fF
C1331 vdd inv_3/in 0.30fF
C1332 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.75fF
C1333 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# clk 0.06fF
C1334 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.06fF
C1335 cla_0/l sumffo_3/k 0.06fF
C1336 ffo_0/nand_1/b ffo_0/nand_7/a 0.13fF
C1337 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_1/op 0.52fF
C1338 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C1339 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b 0.32fF
C1340 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.31fF
C1341 inv_4/in cla_1/n 0.02fF
C1342 sumffo_3/ffo_0/nand_4/w_0_0# sumffo_3/ffo_0/nand_3/b 0.06fF
C1343 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C1344 cla_1/nand_0/w_0_0# gnd 0.01fF
C1345 sumffo_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C1346 ffipgarr_0/ffi_0/nand_0/w_0_0# vdd 0.10fF
C1347 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# vdd 0.11fF
C1348 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# vdd 0.10fF
C1349 cla_1/inv_0/w_0_6# vdd 0.06fF
C1350 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C1351 sumffo_2/xor_0/w_n3_4# inv_2/op 0.06fF
C1352 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/b 0.31fF
C1353 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# vdd 0.10fF
C1354 ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd 0.30fF
C1355 sumffo_0/k vdd 0.31fF
C1356 vdd sumffo_3/ffo_0/inv_0/op 0.17fF
C1357 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C1358 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# vdd 0.10fF
C1359 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.06fF
C1360 y2in clk 0.70fF
C1361 vdd nor_4/a 0.15fF
C1362 vdd sumffo_3/ffo_0/inv_0/w_0_6# 0.06fF
C1363 clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.13fF
C1364 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# vdd 0.10fF
C1365 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.04fF
C1366 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C1367 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d 0.04fF
C1368 sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# 0.02fF
C1369 cla_2/l cla_2/p1 0.02fF
C1370 clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.13fF
C1371 ffipgarr_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.06fF
C1372 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.06fF
C1373 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.06fF
C1374 nand_1/b inv_1/in 0.13fF
C1375 sumffo_3/ffo_0/d sumffo_3/ffo_0/inv_0/w_0_6# 0.06fF
C1376 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/q 0.20fF
C1377 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/w_0_0# 0.06fF
C1378 vdd sumffo_3/ffo_0/nand_7/a 0.30fF
C1379 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C1380 sumffo_2/xor_0/w_n3_4# sumffo_2/k 0.06fF
C1381 sumffo_2/ffo_0/nand_7/a gnd 0.03fF
C1382 ffipgarr_0/ffipg_3/ffi_0/q sumffo_3/k 0.07fF
C1383 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# vdd 0.10fF
C1384 x2in vdd 0.04fF
C1385 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# sumffo_3/k 0.02fF
C1386 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# gnd 0.01fF
C1387 cla_0/n inv_3/w_0_6# 0.00fF
C1388 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/d 0.06fF
C1389 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# vdd 0.93fF
C1390 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C1391 nor_0/a sumffo_1/k 0.06fF
C1392 clk ffo_0/nand_6/a 0.13fF
C1393 ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd 0.03fF
C1394 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.31fF
C1395 ffipgarr_0/ffipg_0/ffi_0/nand_1/b gnd 0.26fF
C1396 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.06fF
C1397 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C1398 sumffo_1/ffo_0/nand_6/a sumffo_1/sbar 0.00fF
C1399 sumffo_2/sbar z3o 0.32fF
C1400 cla_2/g1 gnd 0.27fF
C1401 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# vdd 0.06fF
C1402 vdd gnd 7.10fF
C1403 ffipgarr_0/ffipg_3/ffi_0/inv_1/op gnd 0.22fF
C1404 vdd ffo_0/nand_1/b 0.31fF
C1405 gnd sumffo_1/ffo_0/nand_1/b 0.26fF
C1406 sumffo_0/ffo_0/inv_0/w_0_6# vdd 0.06fF
C1407 ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd 0.03fF
C1408 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/q 0.20fF
C1409 ffipgarr_0/ffipg_2/ffi_0/q gnd 2.62fF
C1410 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.00fF
C1411 gnd sumffo_3/ffo_0/d 0.37fF
C1412 cla_2/g0 cla_2/nor_1/w_0_0# 0.06fF
C1413 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.00fF
C1414 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.04fF
C1415 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C1416 cla_0/nor_1/w_0_0# vdd 0.31fF
C1417 cla_1/g0 gnd 0.76fF
C1418 cla_1/p0 cla_2/p0 0.24fF
C1419 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1420 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.00fF
C1421 ffipgarr_0/ffipg_0/ffi_0/qbar gnd 0.34fF
C1422 cla_2/g1 cla_2/nand_0/w_0_0# 0.06fF
C1423 cla_2/nand_0/w_0_0# vdd 0.10fF
C1424 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# vdd 0.93fF
C1425 ffipgarr_0/ffipg_3/ffi_1/nand_3/b gnd 0.35fF
C1426 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# vdd 0.10fF
C1427 ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd 0.03fF
C1428 ffipgarr_0/ffipg_0/ffi_1/q vdd 1.35fF
C1429 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.32fF
C1430 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.06fF
C1431 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C1432 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C1433 nor_4/b inv_9/in 0.16fF
C1434 gnd ffo_0/nand_3/a 0.14fF
C1435 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/d 0.06fF
C1436 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.04fF
C1437 cla_0/g0 nand_2/b 1.01fF
C1438 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C1439 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# vdd 0.10fF
C1440 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C1441 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# vdd 0.10fF
C1442 cla_0/n inv_5/in 0.13fF
C1443 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk 0.07fF
C1444 ffo_0/nand_7/w_0_0# ffo_0/nand_7/a 0.06fF
C1445 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b 0.13fF
C1446 clk sumffo_2/ffo_0/nand_3/b 0.33fF
C1447 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C1448 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.04fF
C1449 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.06fF
C1450 inv_4/op sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C1451 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C1452 sumffo_2/ffo_0/nand_6/a vdd 0.30fF
C1453 ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd 0.34fF
C1454 vdd sumffo_1/ffo_0/nand_3/w_0_0# 0.11fF
C1455 sumffo_0/xor_0/w_n3_4# vdd 0.12fF
C1456 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op sumffo_3/k 0.52fF
C1457 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# vdd 0.06fF
C1458 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C1459 cla_1/nor_1/w_0_0# vdd 0.31fF
C1460 ffipgarr_0/ffi_0/nand_7/a nand_1/b 0.00fF
C1461 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/qbar 0.00fF
C1462 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C1463 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.31fF
C1464 inv_8/in nor_4/b 0.04fF
C1465 inv_2/in inv_2/op 0.04fF
C1466 vdd sumffo_1/ffo_0/nand_5/w_0_0# 0.10fF
C1467 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.31fF
C1468 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# vdd 0.06fF
C1469 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_1/b 0.04fF
C1470 sumffo_2/xor_0/inv_0/w_0_6# vdd 0.09fF
C1471 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_1/w_0_6# 0.03fF
C1472 ffipgarr_0/ffipg_3/ffi_1/qbar vdd 0.33fF
C1473 ffipgarr_0/ffipg_3/ffi_1/inv_1/op gnd 0.22fF
C1474 ffipgarr_0/ffi_0/nand_1/b gnd 0.26fF
C1475 cla_0/nor_1/a_13_6# gnd 0.01fF
C1476 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.06fF
C1477 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C1478 nand_1/b sumffo_1/k 0.02fF
C1479 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.00fF
C1480 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# vdd 0.10fF
C1481 vdd sumffo_3/ffo_0/nand_4/w_0_0# 0.10fF
C1482 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C1483 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# vdd 0.06fF
C1484 vdd sumffo_1/ffo_0/d 0.04fF
C1485 ffipgarr_0/ffi_0/nand_3/a vdd 0.30fF
C1486 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# clk 0.06fF
C1487 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.04fF
C1488 cla_0/l sumffo_2/ffo_0/nand_2/w_0_0# 0.17fF
C1489 inv_4/op nor_2/w_0_0# 0.03fF
C1490 clk sumffo_1/ffo_0/nand_0/b 0.04fF
C1491 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C1492 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C1493 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.03fF
C1494 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C1495 ffipgarr_0/ffi_0/nand_6/w_0_0# vdd 0.10fF
C1496 x3in ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C1497 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.04fF
C1498 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# vdd 0.11fF
C1499 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# vdd 0.10fF
C1500 vdd inv_3/w_0_6# 0.15fF
C1501 gnd inv_1/in 0.22fF
C1502 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.06fF
C1503 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# vdd 0.10fF
C1504 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar 0.32fF
C1505 ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd 0.35fF
C1506 x1in ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.04fF
C1507 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.04fF
C1508 sumffo_2/ffo_0/nand_3/b cla_0/n 0.19fF
C1509 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/qbar 0.04fF
C1510 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.13fF
C1511 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C1512 ffipgarr_0/ffipg_2/ffi_1/q gnd 0.93fF
C1513 ffipgarr_0/ffipg_1/ffi_1/q gnd 0.93fF
C1514 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk 0.07fF
C1515 cla_1/inv_0/in cla_2/p0 0.02fF
C1516 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C1517 nand_1/b inv_1/w_0_6# 0.06fF
C1518 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/inv_0/op 0.06fF
C1519 ffipgarr_0/ffi_0/nand_5/w_0_0# vdd 0.10fF
C1520 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C1521 y2in vdd 0.04fF
C1522 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C1523 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# gnd 0.00fF
C1524 clk ffipgarr_0/ffi_0/inv_1/op 0.10fF
C1525 ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd 0.30fF
C1526 ffipgarr_0/ffipg_0/ffi_1/nand_1/a clk 0.13fF
C1527 vdd nor_0/w_0_0# 0.15fF
C1528 vdd sumffo_2/xor_0/inv_1/op 0.15fF
C1529 sumffo_0/ffo_0/nand_2/w_0_0# vdd 0.10fF
C1530 ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd 0.30fF
C1531 vdd ffo_0/nand_7/w_0_0# 0.12fF
C1532 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C1533 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b 0.13fF
C1534 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_3/b 0.04fF
C1535 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.04fF
C1536 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C1537 ffipgarr_0/ffipg_2/ffi_1/inv_0/op clk 0.32fF
C1538 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.04fF
C1539 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.06fF
C1540 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.06fF
C1541 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C1542 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/ffi_0/inv_0/w_0_6# 0.03fF
C1543 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.04fF
C1544 cla_2/inv_0/in cla_2/g1 0.04fF
C1545 cla_2/inv_0/in vdd 0.05fF
C1546 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.04fF
C1547 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C1548 x3in ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.04fF
C1549 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.31fF
C1550 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C1551 cla_0/g0 ffipgarr_0/ffipg_0/ffi_0/q 1.40fF
C1552 nand_2/b cla_1/l 0.35fF
C1553 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/ffo_0/nand_6/a 0.06fF
C1554 sumffo_1/sbar sumffo_1/ffo_0/nand_7/w_0_0# 0.06fF
C1555 sumffo_1/ffo_0/nand_6/w_0_0# z2o 0.06fF
C1556 vdd inv_5/in 0.30fF
C1557 inv_2/in nor_1/w_0_0# 0.11fF
C1558 vdd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C1559 vdd sumffo_1/xor_0/w_n3_4# 0.12fF
C1560 ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd 0.39fF
C1561 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.06fF
C1562 vdd ffo_0/nand_6/a 0.30fF
C1563 sumffo_3/k sumffo_3/xor_0/inv_1/op 0.06fF
C1564 gnd sumffo_1/ffo_0/nand_6/a 0.03fF
C1565 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/nand_0/b 0.06fF
C1566 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.00fF
C1567 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a 0.13fF
C1568 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.45fF
C1569 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1570 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op 0.06fF
C1571 ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1572 clk ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.32fF
C1573 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C1574 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C1575 cla_2/g0 cla_1/n 0.13fF
C1576 gnd ffo_0/nand_2/w_0_0# 0.00fF
C1577 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# nand_1/b 0.04fF
C1578 ffipgarr_0/ffipg_1/ffi_1/qbar gnd 0.34fF
C1579 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.31fF
C1580 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.06fF
C1581 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C1582 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C1583 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C1584 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.04fF
C1585 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C1586 vdd nor_2/w_0_0# 0.15fF
C1587 gnd sumffo_3/ffo_0/nand_0/b 0.38fF
C1588 ffipgarr_0/ffi_0/nand_7/a gnd 0.03fF
C1589 ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd 0.22fF
C1590 ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd 0.35fF
C1591 ffipgarr_0/ffipg_0/ffi_0/inv_0/op clk 0.32fF
C1592 cla_1/p0 vdd 0.44fF
C1593 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op nand_1/b 0.04fF
C1594 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.31fF
C1595 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# vdd 0.10fF
C1596 ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd 0.03fF
C1597 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# vdd 0.06fF
C1598 sumffo_2/xor_0/inv_0/op gnd 0.17fF
C1599 sumffo_0/ffo_0/nand_7/a z1o 0.00fF
C1600 nor_4/a inv_9/in 0.02fF
C1601 gnd ffo_0/nand_1/a 0.03fF
C1602 ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd 0.34fF
C1603 gnd sumffo_1/k 0.35fF
C1604 ffipgarr_0/ffipg_1/ffi_0/q vdd 0.38fF
C1605 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1606 ffo_0/d ffo_0/nand_0/b 0.40fF
C1607 clk sumffo_0/ffo_0/nand_1/b 0.45fF
C1608 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C1609 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C1610 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.45fF
C1611 cla_1/g0 cla_1/p0 1.76fF
C1612 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.04fF
C1613 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.06fF
C1614 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.04fF
C1615 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C1616 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.13fF
C1617 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C1618 cla_0/l cla_1/n 0.18fF
C1619 gnd nor_1/b 0.10fF
C1620 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C1621 sumffo_2/ffo_0/nand_3/b vdd 0.39fF
C1622 cla_2/g0 cla_2/p1 0.30fF
C1623 ffipgarr_0/ffipg_3/ffi_1/nand_6/a gnd 0.03fF
C1624 ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd 1.63fF
C1625 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q 0.29fF
C1626 ffo_0/qbar couto 0.32fF
C1627 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C1628 ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd 0.34fF
C1629 cla_0/g0 nor_0/a 1.58fF
C1630 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.06fF
C1631 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.04fF
C1632 cla_2/l cla_0/l 0.40fF
C1633 sumffo_0/sbar vdd 0.28fF
C1634 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# vdd 0.10fF
C1635 sumffo_2/ffo_0/nand_0/w_0_0# cla_0/n 0.04fF
C1636 vdd sumffo_3/ffo_0/nand_2/w_0_0# 0.10fF
C1637 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C1638 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# vdd 0.10fF
C1639 cla_0/nand_0/w_0_0# vdd 0.10fF
C1640 ffipgarr_0/ffi_0/inv_0/op cinin 0.04fF
C1641 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.04fF
C1642 x3in clk 0.70fF
C1643 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C1644 ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd 0.03fF
C1645 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# sumffo_0/k 0.45fF
C1646 gnd inv_1/w_0_6# 0.01fF
C1647 sumffo_3/ffo_0/nand_7/a z4o 0.00fF
C1648 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.06fF
C1649 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# vdd 0.10fF
C1650 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.31fF
C1651 cla_1/n nor_2/b 0.37fF
C1652 sumffo_2/xor_0/a_10_10# vdd 0.93fF
C1653 gnd inv_9/in 0.24fF
C1654 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C1655 vdd sumffo_1/ffo_0/nand_0/b 0.15fF
C1656 sumffo_0/ffo_0/nand_0/b gnd 0.38fF
C1657 ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd 0.39fF
C1658 gnd sumffo_3/k 0.35fF
C1659 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C1660 x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.04fF
C1661 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# vdd 0.10fF
C1662 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/d 0.06fF
C1663 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# gnd 0.00fF
C1664 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.33fF
C1665 cla_0/nand_0/w_0_0# cla_1/g0 0.06fF
C1666 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k 0.06fF
C1667 vdd ffo_0/nand_3/w_0_0# 0.11fF
C1668 sumffo_0/xor_0/inv_0/op vdd 0.15fF
C1669 ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd 0.34fF
C1670 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# vdd 0.06fF
C1671 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C1672 inv_0/op gnd 0.10fF
C1673 inv_4/op sumffo_3/xor_0/inv_0/op 0.20fF
C1674 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/xor_0/inv_0/op 0.03fF
C1675 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.13fF
C1676 y1in gnd 0.19fF
C1677 cla_0/l cla_1/nand_0/a_13_n26# 0.01fF
C1678 ffipgarr_0/ffipg_2/ffi_1/nand_1/a clk 0.13fF
C1679 ffipgarr_0/ffipg_1/ffi_0/nand_3/a clk 0.13fF
C1680 ffo_0/nand_6/w_0_0# ffo_0/qbar 0.04fF
C1681 gnd z4o 0.52fF
C1682 inv_4/in nor_2/b 0.16fF
C1683 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# sumffo_3/k 0.45fF
C1684 ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd 0.10fF
C1685 ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd 1.63fF
C1686 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C1687 cla_1/inv_0/in vdd 0.05fF
C1688 gnd inv_8/in 0.13fF
C1689 cla_2/nand_0/a_13_n26# gnd 0.01fF
C1690 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/qbar 0.00fF
C1691 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.06fF
C1692 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.06fF
C1693 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C1694 cla_2/p1 cla_2/nor_0/w_0_0# 0.06fF
C1695 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# vdd 0.10fF
C1696 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C1697 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.17fF
C1698 ffipgarr_0/ffi_0/inv_1/op vdd 1.67fF
C1699 ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd 0.15fF
C1700 clk cla_0/n 0.12fF
C1701 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# vdd 0.10fF
C1702 x1in gnd 0.19fF
C1703 ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd 0.30fF
C1704 cla_1/g0 cla_1/inv_0/in 0.16fF
C1705 vdd ffo_0/inv_0/op 0.17fF
C1706 cla_1/p0 ffipgarr_0/ffipg_1/ffi_1/q 0.22fF
C1707 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.06fF
C1708 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.06fF
C1709 ffo_0/nand_3/w_0_0# ffo_0/nand_3/a 0.06fF
C1710 sumffo_0/ffo_0/inv_0/op gnd 0.10fF
C1711 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.06fF
C1712 ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd 0.17fF
C1713 ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd 0.03fF
C1714 nand_2/b cla_0/nand_0/a_13_n26# 0.00fF
C1715 cla_0/g0 cla_0/inv_0/in 0.16fF
C1716 cla_0/g0 nand_1/b 0.05fF
C1717 clk sumffo_0/ffo_0/d 0.25fF
C1718 nor_0/b inv_0/in 0.16fF
C1719 sumffo_2/ffo_0/nand_2/w_0_0# sumffo_2/ffo_0/nand_3/a 0.04fF
C1720 ffipgarr_0/ffipg_3/ffi_0/q cla_2/p1 0.03fF
C1721 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/nand_7/a 0.04fF
C1722 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.31fF
C1723 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.13fF
C1724 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.00fF
C1725 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.04fF
C1726 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_1/q 0.73fF
C1727 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/inv_0/w_0_6# 0.03fF
C1728 ffipgarr_0/ffipg_3/ffi_1/q vdd 1.35fF
C1729 y3in ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.01fF
C1730 cla_2/inv_0/op vdd 0.17fF
C1731 cla_2/g1 cla_2/inv_0/op 0.35fF
C1732 ffipgarr_0/ffipg_2/ffi_0/inv_0/op clk 0.32fF
C1733 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C1734 inv_7/op inv_8/w_0_6# 0.06fF
C1735 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_1/op 0.52fF
C1736 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C1737 gnd sumffo_1/ffo_0/nand_3/b 0.35fF
C1738 clk sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C1739 x4in ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C1740 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# clk 0.06fF
C1741 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op gnd 0.17fF
C1742 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C1743 cla_0/g0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C1744 vdd z2o 0.28fF
C1745 z1o gnd 0.52fF
C1746 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op vdd 0.15fF
C1747 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.04fF
C1748 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C1749 sumffo_3/ffo_0/nand_1/w_0_0# sumffo_3/ffo_0/nand_3/b 0.04fF
C1750 sumffo_2/ffo_0/inv_0/op vdd 0.17fF
C1751 ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd 0.17fF
C1752 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/ffo_0/nand_7/a 0.06fF
C1753 sumffo_2/sbar gnd 0.34fF
C1754 sumffo_2/ffo_0/nand_0/w_0_0# vdd 0.10fF
C1755 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.33fF
C1756 ffipgarr_0/ffipg_2/ffi_0/qbar gnd 0.34fF
C1757 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# cla_2/g0 0.04fF
C1758 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1759 nor_3/w_0_0# cla_2/n 0.06fF
C1760 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C1761 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C1762 vdd sumffo_3/sbar 0.28fF
C1763 ffipgarr_0/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C1764 ffipgarr_0/ffipg_3/ffi_0/nand_1/b gnd 0.26fF
C1765 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.06fF
C1766 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C1767 gnd ffo_0/nand_3/b 0.35fF
C1768 sumffo_1/xor_0/w_n3_4# sumffo_1/k 0.06fF
C1769 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C1770 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.06fF
C1771 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.06fF
C1772 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_1/b 0.45fF
C1773 ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd 0.17fF
C1774 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# x2in 0.06fF
C1775 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C1776 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C1777 cla_2/l inv_5/w_0_6# 0.29fF
C1778 vdd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C1779 ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd 0.34fF
C1780 ffo_0/nand_3/b ffo_0/nand_1/b 0.32fF
C1781 vdd sumffo_3/xor_0/inv_0/op 0.15fF
C1782 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op nand_1/b 0.04fF
C1783 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/b 0.31fF
C1784 sumffo_0/ffo_0/nand_1/b vdd 0.31fF
C1785 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C1786 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C1787 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.31fF
C1788 nand_2/b inv_2/op 0.10fF
C1789 sumffo_2/ffo_0/nand_1/w_0_0# cla_0/n 0.13fF
C1790 vdd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C1791 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C1792 ffipgarr_0/ffipg_3/ffi_0/qbar gnd 0.34fF
C1793 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.00fF
C1794 inv_7/op vdd 0.15fF
C1795 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# x1in 0.06fF
C1796 cla_2/nor_1/w_0_0# gnd 0.01fF
C1797 cla_2/l nor_3/b 0.27fF
C1798 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op 0.06fF
C1799 ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd 0.39fF
C1800 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_3/b 0.00fF
C1801 cla_1/p0 sumffo_1/k 0.05fF
C1802 inv_9/in Gnd 0.23fF
C1803 nor_4/w_0_0# Gnd 1.81fF
C1804 nor_4/b Gnd 1.06fF
C1805 inv_8/in Gnd 0.22fF
C1806 inv_8/w_0_6# Gnd 1.40fF
C1807 inv_7/in Gnd 0.22fF
C1808 inv_7/w_0_6# Gnd 1.40fF
C1809 nor_4/a Gnd 0.27fF
C1810 inv_5/in Gnd 0.22fF
C1811 inv_5/w_0_6# Gnd 1.40fF
C1812 nor_3/b Gnd 0.92fF
C1813 cla_2/n Gnd 0.32fF
C1814 inv_6/in Gnd 0.23fF
C1815 nor_3/w_0_0# Gnd 1.81fF
C1816 nor_2/b Gnd 0.92fF
C1817 cla_1/n Gnd 0.20fF
C1818 inv_4/in Gnd 0.23fF
C1819 nor_2/w_0_0# Gnd 1.81fF
C1820 inv_3/in Gnd 0.22fF
C1821 inv_3/w_0_6# Gnd 1.40fF
C1822 inv_2/op Gnd 1.94fF
C1823 inv_2/in Gnd 0.23fF
C1824 nor_1/w_0_0# Gnd 1.81fF
C1825 nor_1/b Gnd 0.85fF
C1826 inv_1/in Gnd 0.22fF
C1827 inv_1/w_0_6# Gnd 1.40fF
C1828 inv_0/in Gnd 0.23fF
C1829 nor_0/w_0_0# Gnd 1.81fF
C1830 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1831 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1832 ffo_0/nand_7/a Gnd 0.30fF
C1833 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1834 ffo_0/qbar Gnd 0.42fF
C1835 ffo_0/nand_6/a Gnd 0.30fF
C1836 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1837 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1838 ffo_0/nand_3/b Gnd 0.43fF
C1839 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1840 ffo_0/nand_3/a Gnd 0.30fF
C1841 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1842 ffo_0/nand_0/b Gnd 0.63fF
C1843 ffo_0/d Gnd 0.60fF
C1844 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1845 ffo_0/inv_0/op Gnd 0.26fF
C1846 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1847 ffo_0/nand_1/a Gnd 0.30fF
C1848 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1849 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1850 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1851 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1852 inv_4/op Gnd 1.54fF
C1853 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1854 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1855 sumffo_3/k Gnd 3.28fF
C1856 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1857 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1858 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1859 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1860 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1861 sumffo_3/sbar Gnd 0.43fF
C1862 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1863 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1864 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1865 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1866 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1867 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1868 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1869 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1870 sumffo_3/ffo_0/d Gnd 0.64fF
C1871 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1872 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1873 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1874 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1875 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1876 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1877 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1878 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1879 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1880 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1881 sumffo_1/k Gnd 2.61fF
C1882 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1883 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1884 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1885 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1886 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1887 sumffo_1/sbar Gnd 0.43fF
C1888 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1889 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1890 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1891 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1892 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1893 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1894 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1895 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1896 sumffo_1/ffo_0/d Gnd 0.64fF
C1897 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1898 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1899 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1900 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1901 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1902 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1903 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1904 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1905 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1906 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1907 sumffo_2/k Gnd 1.72fF
C1908 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1909 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1910 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1911 gnd Gnd 46.05fF
C1912 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1913 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1914 sumffo_2/sbar Gnd 0.43fF
C1915 vdd Gnd 27.12fF
C1916 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1917 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1918 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1919 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1920 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1921 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1922 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1923 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1924 sumffo_2/ffo_0/d Gnd 0.64fF
C1925 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1926 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1927 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1928 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1929 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1930 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1931 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1932 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1933 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1934 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1935 sumffo_0/k Gnd 3.08fF
C1936 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1937 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1938 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1939 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1940 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1941 sumffo_0/sbar Gnd 0.43fF
C1942 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1943 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1944 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1945 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1946 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1947 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1948 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1949 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1950 sumffo_0/ffo_0/d Gnd 0.64fF
C1951 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1952 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1953 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1954 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1955 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1956 cla_2/p1 Gnd 1.08fF
C1957 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1958 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1959 cla_2/inv_0/in Gnd 0.27fF
C1960 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1961 cla_2/g1 Gnd 0.58fF
C1962 cla_2/inv_0/op Gnd 0.26fF
C1963 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1964 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1965 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1966 ffipgarr_0/ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1967 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1968 ffipgarr_0/ffipg_3/ffi_1/qbar Gnd 0.42fF
C1969 ffipgarr_0/ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1970 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1971 ffipgarr_0/ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1972 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1973 ffipgarr_0/ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1974 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1975 ffipgarr_0/ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1976 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1977 x4in Gnd 0.52fF
C1978 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1979 ffipgarr_0/ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1980 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1981 ffipgarr_0/ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1982 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1983 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1984 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1985 ffipgarr_0/ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1986 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1987 ffipgarr_0/ffipg_3/ffi_0/qbar Gnd 0.42fF
C1988 ffipgarr_0/ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1989 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1990 ffipgarr_0/ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1991 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1992 ffipgarr_0/ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1993 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1994 ffipgarr_0/ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1995 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1996 y4in Gnd 0.52fF
C1997 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1998 ffipgarr_0/ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1999 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2000 ffipgarr_0/ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C2001 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2002 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2003 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2004 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2005 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2006 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2007 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2008 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2009 ffipgarr_0/ffipg_3/ffi_0/q Gnd 2.68fF
C2010 ffipgarr_0/ffipg_3/ffi_1/q Gnd 2.93fF
C2011 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2012 ffipgarr_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2013 ffipgarr_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2014 ffipgarr_0/ffi_0/nand_7/a Gnd 0.30fF
C2015 ffipgarr_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2016 nor_0/b Gnd 1.09fF
C2017 ffipgarr_0/ffi_0/nand_6/a Gnd 0.30fF
C2018 ffipgarr_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2019 ffipgarr_0/ffi_0/inv_1/op Gnd 0.89fF
C2020 ffipgarr_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2021 ffipgarr_0/ffi_0/nand_3/b Gnd 0.43fF
C2022 ffipgarr_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2023 ffipgarr_0/ffi_0/nand_3/a Gnd 0.30fF
C2024 ffipgarr_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2025 clk Gnd 17.25fF
C2026 cinin Gnd 0.52fF
C2027 ffipgarr_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2028 ffipgarr_0/ffi_0/inv_0/op Gnd 0.26fF
C2029 ffipgarr_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2030 ffipgarr_0/ffi_0/nand_1/a Gnd 0.30fF
C2031 ffipgarr_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2032 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2033 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2034 ffipgarr_0/ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C2035 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2036 ffipgarr_0/ffipg_2/ffi_1/qbar Gnd 0.42fF
C2037 ffipgarr_0/ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C2038 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2039 ffipgarr_0/ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C2040 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2041 ffipgarr_0/ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C2042 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2043 ffipgarr_0/ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C2044 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2045 x3in Gnd 0.52fF
C2046 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2047 ffipgarr_0/ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C2048 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2049 ffipgarr_0/ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C2050 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2051 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2052 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2053 ffipgarr_0/ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C2054 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2055 ffipgarr_0/ffipg_2/ffi_0/qbar Gnd 0.42fF
C2056 ffipgarr_0/ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C2057 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2058 ffipgarr_0/ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C2059 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2060 ffipgarr_0/ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C2061 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2062 ffipgarr_0/ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C2063 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2064 y3in Gnd 0.52fF
C2065 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2066 ffipgarr_0/ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C2067 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2068 ffipgarr_0/ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C2069 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2070 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2071 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2072 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2073 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2074 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2075 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2076 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2077 ffipgarr_0/ffipg_2/ffi_0/q Gnd 2.68fF
C2078 ffipgarr_0/ffipg_2/ffi_1/q Gnd 2.93fF
C2079 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2080 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2081 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2082 ffipgarr_0/ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C2083 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2084 ffipgarr_0/ffipg_1/ffi_1/qbar Gnd 0.42fF
C2085 ffipgarr_0/ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C2086 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2087 ffipgarr_0/ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C2088 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2089 ffipgarr_0/ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C2090 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2091 ffipgarr_0/ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C2092 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2093 x2in Gnd 0.52fF
C2094 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2095 ffipgarr_0/ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C2096 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2097 ffipgarr_0/ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C2098 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2099 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2100 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2101 ffipgarr_0/ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C2102 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2103 ffipgarr_0/ffipg_1/ffi_0/qbar Gnd 0.42fF
C2104 ffipgarr_0/ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C2105 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2106 ffipgarr_0/ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C2107 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2108 ffipgarr_0/ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C2109 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2110 ffipgarr_0/ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C2111 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2112 y2in Gnd 0.43fF
C2113 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2114 ffipgarr_0/ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C2115 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2116 ffipgarr_0/ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C2117 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2118 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2119 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2120 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2121 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2122 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2123 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2124 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2125 ffipgarr_0/ffipg_1/ffi_0/q Gnd 2.68fF
C2126 ffipgarr_0/ffipg_1/ffi_1/q Gnd 2.93fF
C2127 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2128 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2129 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2130 ffipgarr_0/ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C2131 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2132 ffipgarr_0/ffipg_0/ffi_1/qbar Gnd 0.42fF
C2133 ffipgarr_0/ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C2134 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2135 ffipgarr_0/ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C2136 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2137 ffipgarr_0/ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C2138 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2139 ffipgarr_0/ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C2140 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2141 x1in Gnd 0.42fF
C2142 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2143 ffipgarr_0/ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C2144 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2145 ffipgarr_0/ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C2146 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2147 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2148 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2149 ffipgarr_0/ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C2150 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2151 ffipgarr_0/ffipg_0/ffi_0/qbar Gnd 0.42fF
C2152 ffipgarr_0/ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C2153 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2154 ffipgarr_0/ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C2155 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2156 ffipgarr_0/ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C2157 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2158 ffipgarr_0/ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C2159 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2160 y1in Gnd 0.52fF
C2161 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2162 ffipgarr_0/ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C2163 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2164 ffipgarr_0/ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C2165 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2166 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2167 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2168 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2169 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2170 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2171 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2172 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2173 ffipgarr_0/ffipg_0/ffi_0/q Gnd 2.68fF
C2174 ffipgarr_0/ffipg_0/ffi_1/q Gnd 2.93fF
C2175 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2176 cla_1/nor_1/w_0_0# Gnd 1.23fF
C2177 cla_1/l Gnd 0.31fF
C2178 cla_1/nor_0/w_0_0# Gnd 1.23fF
C2179 cla_1/inv_0/in Gnd 0.27fF
C2180 cla_1/inv_0/w_0_6# Gnd 0.58fF
C2181 cla_1/inv_0/op Gnd 0.26fF
C2182 cla_1/nand_0/w_0_0# Gnd 0.82fF
C2183 inv_7/op Gnd 0.30fF
C2184 nand_5/a Gnd 0.16fF
C2185 cla_0/nor_1/w_0_0# Gnd 1.23fF
C2186 cla_0/l Gnd 7.05fF
C2187 cla_0/nor_0/w_0_0# Gnd 1.23fF
C2188 cla_0/inv_0/in Gnd 0.27fF
C2189 cla_0/inv_0/w_0_6# Gnd 0.58fF
C2190 cla_1/g0 Gnd 2.32fF
C2191 cla_0/inv_0/op Gnd 0.26fF
C2192 cla_0/nand_0/w_0_0# Gnd 0.82fF
C2193 cla_2/l Gnd 1.05fF
C2194 nand_2/b Gnd 0.27fF
C2195 inv_0/op Gnd 0.26fF
C2196 nand_0/w_0_0# Gnd 0.82fF
