* SPICE3 file created from tspc.ext - technology: scmos

.option scale=0.01u

M1000 clk clk gnd Gnd nfet w=54 l=18
+  ad=2430 pd=198 as=17010 ps=1116
M1001 clk clk vdd inv_0/w_0_6# pfet w=108 l=18
+  ad=4860 pd=306 as=21870 ps=1332
M1002 a_n69_1# d gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1003 d a_13_35# vdd w_0_29# pfet w=126 l=18
+  ad=34020 pd=1044 as=0 ps=0
M1004 a_13_1# d gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1005 d clk a_n35_1# Gnd nfet w=108 l=18
+  ad=13608 pd=684 as=5832 ps=324
M1006 a_13_35# d vdd w_0_29# pfet w=126 l=18
+  ad=17010 pd=522 as=0 ps=0
M1007 a_13_35# clk a_13_1# Gnd nfet w=108 l=18
+  ad=6804 pd=342 as=0 ps=0
M1008 a_n35_1# a_n69_35# gnd Gnd nfet w=108 l=18
+  ad=0 pd=0 as=0 ps=0
M1009 a_n69_35# d vdd w_n82_29# pfet w=126 l=18
+  ad=17010 pd=522 as=0 ps=0
M1010 a_47_1# a_13_35# gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1011 a_n69_35# clk a_n69_1# Gnd nfet w=108 l=18
+  ad=6804 pd=342 as=0 ps=0
M1012 d clk a_47_1# Gnd nfet w=108 l=18
+  ad=0 pd=0 as=0 ps=0
M1013 d a_n69_35# vdd w_n82_29# pfet w=126 l=18
+  ad=0 pd=0 as=0 ps=0
C0 d clk 0.98fF
C1 d inv_0/w_0_6# 0.13fF
C2 vdd a_n69_35# 0.03fF
C3 inv_0/w_0_6# clk 0.31fF
C4 d vdd 0.13fF
C5 w_n82_29# a_n69_35# 0.10fF
C6 a_13_35# clk 0.46fF
C7 clk a_n35_1# 0.01fF
C8 clk vdd 0.17fF
C9 inv_0/w_0_6# vdd 0.06fF
C10 w_n82_29# d 0.10fF
C11 a_13_35# vdd 0.03fF
C12 w_0_29# d 0.10fF
C13 gnd a_n69_35# 0.03fF
C14 a_n69_1# clk 0.01fF
C15 w_n82_29# vdd 0.14fF
C16 a_13_35# w_0_29# 0.10fF
C17 d gnd 0.07fF
C18 w_0_29# vdd 0.14fF
C19 gnd clk 0.47fF
C20 clk a_n69_35# 0.54fF
C21 a_13_35# gnd 0.03fF
C22 d Gnd 0.89fF
C23 w_0_29# Gnd 0.39fF
C24 w_n82_29# Gnd 0.39fF
C25 gnd Gnd 0.29fF
C26 clk Gnd 2.64fF
C27 vdd Gnd 0.18fF
C28 inv_0/w_0_6# Gnd 0.58fF
