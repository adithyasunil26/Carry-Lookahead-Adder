* SPICE3 file created from ffo.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=540 ps=316
M1001 vdd nand_1/b nand_3/b nand_1/w_0_0# pfet w=12 l=2
+  ad=1080 pd=612 as=96 ps=40
M1002 nand_3/b nand_1/a vdd nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 nand_3/b nand_1/b nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd nand_0/b nand_1/a nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_1/a inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_1/a nand_0/b nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_0/b nand_3/a nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 nand_3/a d vdd nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 nand_3/a nand_0/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd nand_3/b nand_1/b nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 nand_1/b nand_3/a vdd nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 nand_1/b nand_3/b nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd clk nand_6/a nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 nand_6/a nand_3/b vdd nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 nand_6/a clk nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd nand_1/b nand_7/a nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 nand_7/a clk vdd nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 nand_7/a nand_1/b nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 nand_6/a_13_n26# nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1025 vdd qbar q nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1026 q nand_6/a vdd nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 q qbar nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1028 nand_7/a_13_n26# nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1029 vdd q qbar nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1030 qbar nand_7/a vdd nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 qbar q nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1032 inv_0/op d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1033 inv_0/op d vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1034 nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1035 nand_0/b clk vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 nand_3/a nand_2/w_0_0# 0.04fF
C1 nand_6/a clk 0.13fF
C2 d vdd 0.04fF
C3 qbar nand_7/a 0.00fF
C4 qbar vdd 0.28fF
C5 gnd clk 0.17fF
C6 inv_0/w_0_6# d 0.06fF
C7 nand_0/w_0_0# nand_1/a 0.04fF
C8 inv_1/w_0_6# clk 0.06fF
C9 gnd nand_6/a 0.03fF
C10 nand_3/b clk 0.33fF
C11 nand_0/w_0_0# nand_0/b 0.06fF
C12 nand_0/b clk 0.04fF
C13 nand_2/w_0_0# vdd 0.10fF
C14 nand_4/w_0_0# vdd 0.10fF
C15 qbar nand_7/w_0_0# 0.04fF
C16 nand_3/a vdd 0.30fF
C17 nand_6/a nand_6/w_0_0# 0.06fF
C18 gnd nand_1/a 0.03fF
C19 nand_3/b gnd 0.35fF
C20 nand_3/b nand_1/a 0.00fF
C21 inv_0/op vdd 0.17fF
C22 nand_3/a nand_3/w_0_0# 0.06fF
C23 gnd nand_0/b 0.38fF
C24 nand_5/w_0_0# nand_1/b 0.06fF
C25 nand_1/a nand_0/b 0.13fF
C26 nand_5/w_0_0# nand_7/a 0.04fF
C27 inv_1/w_0_6# nand_0/b 0.03fF
C28 nand_7/a q 0.31fF
C29 qbar nand_6/a 0.31fF
C30 nand_5/w_0_0# vdd 0.10fF
C31 q vdd 0.28fF
C32 nand_1/a nand_1/w_0_0# 0.06fF
C33 inv_0/w_0_6# inv_0/op 0.03fF
C34 nand_3/b nand_1/w_0_0# 0.04fF
C35 nand_7/a nand_1/b 0.13fF
C36 gnd d 0.16fF
C37 vdd nand_1/b 0.31fF
C38 gnd qbar 0.52fF
C39 nand_7/a vdd 0.30fF
C40 nand_0/b d 0.40fF
C41 nand_4/w_0_0# clk 0.06fF
C42 nand_3/w_0_0# nand_1/b 0.04fF
C43 nand_4/w_0_0# nand_6/a 0.04fF
C44 nand_3/w_0_0# vdd 0.11fF
C45 nand_7/w_0_0# q 0.06fF
C46 qbar nand_6/w_0_0# 0.06fF
C47 inv_0/w_0_6# vdd 0.06fF
C48 nand_0/w_0_0# inv_0/op 0.06fF
C49 nand_5/w_0_0# clk 0.06fF
C50 nand_7/a nand_7/w_0_0# 0.06fF
C51 nand_3/a gnd 0.03fF
C52 nand_7/w_0_0# vdd 0.10fF
C53 q nand_6/a 0.00fF
C54 nand_3/b nand_4/w_0_0# 0.06fF
C55 nand_3/b nand_3/a 0.31fF
C56 gnd inv_0/op 0.10fF
C57 nand_0/b nand_2/w_0_0# 0.06fF
C58 nand_3/a nand_0/b 0.13fF
C59 nand_1/b clk 0.45fF
C60 nand_0/w_0_0# vdd 0.10fF
C61 vdd clk 1.49fF
C62 gnd q 0.34fF
C63 vdd nand_6/a 0.30fF
C64 nand_0/b inv_0/op 0.32fF
C65 d nand_2/w_0_0# 0.06fF
C66 gnd nand_1/b 0.26fF
C67 nand_1/a nand_1/b 0.31fF
C68 gnd nand_7/a 0.03fF
C69 gnd vdd 0.03fF
C70 q nand_6/w_0_0# 0.04fF
C71 d inv_0/op 0.04fF
C72 nand_3/b nand_1/b 0.32fF
C73 nand_1/a vdd 0.30fF
C74 inv_1/w_0_6# vdd 0.06fF
C75 nand_3/b vdd 0.39fF
C76 nand_0/b vdd 0.15fF
C77 nand_1/w_0_0# nand_1/b 0.06fF
C78 qbar q 0.32fF
C79 vdd nand_6/w_0_0# 0.10fF
C80 nand_3/b nand_3/w_0_0# 0.06fF
C81 nand_1/w_0_0# vdd 0.10fF
C82 inv_1/w_0_6# Gnd 0.58fF
C83 inv_0/w_0_6# Gnd 0.58fF
C84 gnd Gnd 1.75fF
C85 nand_7/a Gnd 0.30fF
C86 nand_7/w_0_0# Gnd 0.82fF
C87 q Gnd 0.42fF
C88 vdd Gnd 1.12fF
C89 nand_6/a Gnd 0.30fF
C90 nand_6/w_0_0# Gnd 0.82fF
C91 clk Gnd 1.05fF
C92 nand_5/w_0_0# Gnd 0.82fF
C93 nand_3/b Gnd 0.43fF
C94 nand_4/w_0_0# Gnd 0.82fF
C95 nand_3/a Gnd 0.30fF
C96 nand_3/w_0_0# Gnd 0.82fF
C97 nand_0/b Gnd 0.63fF
C98 d Gnd 0.45fF
C99 nand_2/w_0_0# Gnd 0.82fF
C100 inv_0/op Gnd 0.26fF
C101 nand_0/w_0_0# Gnd 0.82fF
C102 nand_1/a Gnd 0.30fF
C103 nand_1/w_0_0# Gnd 0.82fF
