* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 gnd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 gnd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 gnd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 gnd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 gnd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 gnd cla_0/l cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op gnd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_0/l cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in gnd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=312 pd=138 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 gnd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=168 ps=96
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 gnd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 gnd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 gnd cla_0/l cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op gnd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_0/l cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in gnd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 gnd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_0/l cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 gnd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_0/l cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 gnd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op gnd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in gnd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 gnd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_0/l cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 gnd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_0/l cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin gnd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 gnd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 sumffo_0/xor_0/op cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/op sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k gnd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 sumffo_0/xor_0/op sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op gnd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op ffipg_2/k gnd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 gnd ffipg_2/k sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 sumffo_2/xor_0/op ffipg_2/k sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op gnd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 sumffo_2/xor_0/op sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b gnd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 gnd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 sumffo_1/xor_0/op nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/op sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k gnd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 sumffo_1/xor_0/op sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op gnd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 gnd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 sumffo_3/xor_0/op ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/op sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op gnd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 sumffo_3/xor_0/op sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in gnd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in gnd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in gnd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a gnd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in gnd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n gnd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in gnd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n gnd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in gnd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n gnd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in gnd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a gnd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in gnd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in gnd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 gnd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in gnd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 gnd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in gnd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in gnd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in gnd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 gnd y2in cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 cla_0/l x2in gnd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_0/l y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 gnd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in gnd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in gnd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 gnd y3in cla_0/l ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 cla_0/l x3in gnd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_0/l y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 gnd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in gnd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in gnd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 gnd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in gnd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 gnd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in gnd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in gnd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 cla_2/l inv_5/in 0.05fF
C1 gnd sumffo_3/xor_0/inv_1/op 0.35fF
C2 cla_0/inv_0/in cla_0/l 0.07fF
C3 ffipg_1/pggen_0/xor_0/inv_1/op x2in 0.06fF
C4 sumffo_0/xor_0/op sumffo_0/xor_0/inv_0/op 0.06fF
C5 cin inv_2/in 0.13fF
C6 gnd nor_4/a 0.40fF
C7 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C8 ffipg_1/pggen_0/xor_0/inv_1/op gnd 0.39fF
C9 cin sumffo_1/xor_0/w_n3_4# 0.00fF
C10 gnd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C11 gnd sumffo_1/xor_0/a_10_10# 0.93fF
C12 sumffo_2/xor_0/inv_1/w_0_6# ffipg_2/k 0.23fF
C13 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C14 cla_0/g0 ffipg_1/k 0.06fF
C15 nor_3/w_0_0# gnd 0.14fF
C16 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/op 0.52fF
C17 inv_4/op ffipg_3/k 0.09fF
C18 y4in ffipg_3/k 0.07fF
C19 nor_3/w_0_0# inv_6/in 0.11fF
C20 x1in gnd 1.19fF
C21 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C22 cla_0/l cla_1/nor_1/w_0_0# 0.09fF
C23 x4in gnd 1.24fF
C24 gnd nor_4/w_0_0# 0.15fF
C25 nor_3/b inv_5/w_0_6# 0.17fF
C26 sumffo_0/xor_0/op gnd 0.14fF
C27 nor_0/w_0_0# cin 0.16fF
C28 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/op 0.52fF
C29 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k 0.52fF
C30 gnd nor_3/b 0.33fF
C31 x1in nor_0/a 0.22fF
C32 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C33 nor_3/b inv_6/in 0.16fF
C34 cla_2/g1 gnd 0.65fF
C35 cin sumffo_1/xor_0/op 0.27fF
C36 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k 0.52fF
C37 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.36fF
C38 cla_0/l y3in 0.13fF
C39 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C40 ffipg_0/pggen_0/nor_0/w_0_0# x1in 0.06fF
C41 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.32fF
C42 sumffo_0/xor_0/w_n3_4# ffipg_0/k 0.06fF
C43 gnd cout 0.25fF
C44 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C45 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C46 cla_0/inv_0/op gnd 0.27fF
C47 cin sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C48 sumffo_2/xor_0/inv_0/op cin 0.06fF
C49 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C50 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C51 cla_2/p1 y4in 0.03fF
C52 sumffo_1/xor_0/inv_1/w_0_6# nand_2/b 0.23fF
C53 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C54 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.35fF
C55 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C56 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C57 ffipg_0/pggen_0/xor_0/w_n3_4# y1in 0.06fF
C58 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C59 cla_1/inv_0/in gnd 0.34fF
C60 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C61 cin sumffo_3/xor_0/op 0.16fF
C62 ffipg_0/pggen_0/xor_0/a_10_10# gnd 0.93fF
C63 cla_1/p0 cla_1/l 0.16fF
C64 gnd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C65 cla_1/nand_0/w_0_0# gnd 0.10fF
C66 cla_0/nand_0/w_0_0# cla_0/l 0.06fF
C67 ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C68 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C69 x2in cla_1/p0 0.22fF
C70 cla_0/n inv_5/in 0.13fF
C71 x2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C72 cla_1/p0 gnd 1.12fF
C73 nor_4/a nor_4/w_0_0# 0.07fF
C74 ffipg_1/pggen_0/nor_0/w_0_0# cla_1/p0 0.05fF
C75 ffipg_1/pggen_0/nand_0/w_0_0# gnd 0.10fF
C76 cin sumffo_1/xor_0/inv_0/op 0.06fF
C77 inv_4/op inv_4/in 0.04fF
C78 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C79 cla_1/n cla_1/nand_0/w_0_0# 0.04fF
C80 ffipg_1/pggen_0/xor_0/inv_0/op y2in 0.20fF
C81 gnd sumffo_3/xor_0/inv_0/op 0.32fF
C82 gnd nor_4/b 0.25fF
C83 cla_2/n gnd 0.60fF
C84 cla_1/p0 nor_0/a 0.24fF
C85 ffipg_2/k y3in 0.07fF
C86 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C87 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/k 0.45fF
C88 cla_2/n inv_6/in 0.02fF
C89 inv_6/in nor_4/b 0.04fF
C90 cla_0/l ffipg_3/k 0.10fF
C91 cla_0/l cla_1/inv_0/op 0.35fF
C92 nor_3/w_0_0# nor_3/b 0.06fF
C93 sumffo_2/xor_0/inv_0/op ffipg_2/k 0.20fF
C94 sumffo_2/xor_0/inv_1/w_0_6# gnd 0.06fF
C95 inv_3/in nor_2/b 0.04fF
C96 cla_2/nand_0/a_13_n26# gnd 0.01fF
C97 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C98 cla_0/l nand_2/b 0.06fF
C99 cla_1/p0 ffipg_1/k 0.05fF
C100 cla_2/l cla_2/p1 0.02fF
C101 cin nand_2/b 0.04fF
C102 x1in ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C103 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C104 x4in ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C105 y4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C106 ffipg_0/k y1in 0.07fF
C107 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.39fF
C108 nor_4/w_0_0# cout 0.03fF
C109 cin sumffo_0/xor_0/inv_1/op 0.22fF
C110 cla_2/p0 cla_1/inv_0/in 0.02fF
C111 cla_0/g0 cla_1/p0 0.38fF
C112 gnd nor_2/w_0_0# 0.17fF
C113 cin sumffo_2/xor_0/a_38_n43# 0.01fF
C114 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C115 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/op 0.45fF
C116 cla_0/l y2in 0.13fF
C117 sumffo_2/xor_0/op sumffo_2/xor_0/a_10_10# 0.45fF
C118 cin ffipg_0/k 0.19fF
C119 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C120 cla_0/l cla_2/p1 0.30fF
C121 sumffo_2/xor_0/inv_0/op inv_1/op 0.27fF
C122 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C123 ffipg_0/pggen_0/nand_0/w_0_0# y1in 0.06fF
C124 cla_1/n nor_2/w_0_0# 0.06fF
C125 cla_1/p0 cla_2/p0 0.24fF
C126 cin sumffo_2/xor_0/inv_1/op 0.04fF
C127 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C128 ffipg_3/pggen_0/xor_0/inv_1/op gnd 0.35fF
C129 gnd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C130 cin sumffo_2/xor_0/op 0.28fF
C131 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C132 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/op 0.02fF
C133 gnd inv_2/in 0.47fF
C134 cla_0/inv_0/in gnd 0.34fF
C135 sumffo_2/xor_0/op sumffo_2/xor_0/w_n3_4# 0.02fF
C136 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C137 gnd sumffo_1/xor_0/w_n3_4# 0.12fF
C138 ffipg_2/pggen_0/nand_0/w_0_0# y3in 0.06fF
C139 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# y2in 0.23fF
C140 nand_2/b inv_3/in 0.13fF
C141 nor_4/a nor_4/b 0.42fF
C142 gnd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C143 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_0/op 0.08fF
C144 inv_7/op inv_7/in 0.04fF
C145 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C146 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C147 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.36fF
C148 inv_5/in inv_5/w_0_6# 0.10fF
C149 cla_0/n ffipg_3/k 0.06fF
C150 cla_1/inv_0/op cla_0/n 0.06fF
C151 nor_3/w_0_0# cla_2/n 0.06fF
C152 nor_3/w_0_0# nor_4/b 0.03fF
C153 cla_0/n nor_1/b 0.36fF
C154 cla_2/p1 cla_2/inv_0/in 0.02fF
C155 gnd inv_5/in 0.49fF
C156 cin sumffo_0/xor_0/w_n3_4# 0.06fF
C157 ffipg_2/k nand_2/b 0.06fF
C158 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.15fF
C159 cla_1/nor_1/w_0_0# gnd 0.31fF
C160 nor_0/w_0_0# gnd 0.46fF
C161 inv_7/op cin 0.31fF
C162 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C163 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C164 inv_2/w_0_6# inv_2/in 0.10fF
C165 nor_4/w_0_0# nor_4/b 0.06fF
C166 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C167 cla_0/n nand_2/b 0.06fF
C168 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C169 gnd sumffo_1/xor_0/op 0.14fF
C170 x3in ffipg_2/k 0.46fF
C171 cla_2/n nor_3/b 0.41fF
C172 nor_0/w_0_0# nor_0/a 0.06fF
C173 ffipg_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C174 cla_2/g1 cla_2/n 0.13fF
C175 gnd y3in 1.82fF
C176 ffipg_2/pggen_0/xor_0/a_10_10# gnd 0.93fF
C177 x3in ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C178 cla_0/g0 cla_0/inv_0/in 0.16fF
C179 gnd cinbar 0.16fF
C180 gnd sumffo_0/xor_0/inv_1/w_0_6# 0.07fF
C181 nor_0/w_0_0# inv_0/in 0.11fF
C182 gnd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C183 sumffo_2/xor_0/inv_1/op ffipg_2/k 0.22fF
C184 sumffo_2/xor_0/inv_0/op gnd 0.32fF
C185 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/k 0.01fF
C186 inv_3/w_0_6# nor_2/b 0.03fF
C187 cla_0/n inv_1/in 0.02fF
C188 nor_0/a cinbar 0.32fF
C189 y1in ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C190 cin sumffo_0/xor_0/a_10_10# 0.12fF
C191 nor_0/w_0_0# cla_0/g0 0.06fF
C192 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C193 gnd nor_2/b 0.32fF
C194 inv_8/in cin 0.13fF
C195 inv_0/in cinbar 0.16fF
C196 gnd sumffo_3/xor_0/op 0.14fF
C197 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C198 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C199 ffipg_0/pggen_0/xor_0/w_n3_4# gnd 0.12fF
C200 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C201 ffipg_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C202 cla_1/n nor_2/b 0.39fF
C203 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C204 cla_0/nand_0/w_0_0# gnd 0.10fF
C205 y2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C206 inv_1/op inv_1/in 0.04fF
C207 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C208 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C209 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C210 cla_2/nand_0/w_0_0# gnd 0.18fF
C211 cla_2/l cla_0/l 0.37fF
C212 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C213 gnd sumffo_1/xor_0/inv_0/op 0.32fF
C214 cin sumffo_1/xor_0/inv_1/op 0.04fF
C215 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/inv_0/op 0.08fF
C216 y4in ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C217 x3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C218 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C219 cla_2/p0 y3in 0.03fF
C220 cla_0/l inv_7/in 0.13fF
C221 gnd ffipg_0/pggen_0/nand_0/a_13_n26# 0.01fF
C222 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C223 cin sumffo_2/xor_0/a_10_10# 0.04fF
C224 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C225 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/op 0.45fF
C226 inv_1/op sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C227 inv_7/op inv_7/w_0_6# 0.03fF
C228 gnd ffipg_3/k 0.66fF
C229 cla_1/inv_0/op gnd 0.27fF
C230 nand_2/b inv_3/w_0_6# 0.06fF
C231 gnd nor_1/b 0.35fF
C232 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C233 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C234 cla_1/l nand_2/b 0.31fF
C235 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C236 nor_3/b inv_5/in 0.04fF
C237 sumffo_0/xor_0/inv_0/op ffipg_0/k 0.27fF
C238 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C239 cla_0/l cin 0.33fF
C240 ffipg_2/pggen_0/nor_0/w_0_0# y3in 0.06fF
C241 gnd nand_2/b 1.92fF
C242 cin sumffo_2/xor_0/w_n3_4# 0.00fF
C243 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C244 sumffo_1/xor_0/inv_0/op ffipg_1/k 0.27fF
C245 gnd sumffo_0/xor_0/inv_1/op 0.35fF
C246 ffipg_3/pggen_0/nor_0/w_0_0# ffipg_3/k 0.21fF
C247 inv_8/w_0_6# inv_7/op 0.06fF
C248 x3in gnd 1.24fF
C249 ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/k 0.01fF
C250 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/op 0.52fF
C251 x2in y2in 0.73fF
C252 inv_2/w_0_6# nor_1/b 0.03fF
C253 gnd ffipg_0/k 0.74fF
C254 cla_0/l cla_2/inv_0/in 0.16fF
C255 gnd y2in 1.82fF
C256 nor_1/w_0_0# nor_1/b 0.06fF
C257 ffipg_1/pggen_0/nor_0/w_0_0# y2in 0.06fF
C258 gnd inv_1/in 0.33fF
C259 cla_2/p1 gnd 1.00fF
C260 gnd sumffo_2/xor_0/inv_1/op 0.35fF
C261 gnd sumffo_2/xor_0/op 0.14fF
C262 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C263 cla_0/l cla_2/nor_1/w_0_0# 0.06fF
C264 nand_2/b inv_2/w_0_6# 0.03fF
C265 ffipg_0/k nor_0/a 0.05fF
C266 gnd ffipg_2/pggen_0/nand_0/a_13_n26# 0.01fF
C267 cla_0/inv_0/in cla_1/p0 0.02fF
C268 inv_0/op gnd 0.27fF
C269 ffipg_1/k nand_2/b 0.15fF
C270 cla_0/nand_0/a_13_n26# gnd 0.00fF
C271 gnd ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C272 cla_1/inv_0/w_0_6# gnd 0.06fF
C273 cla_2/l cla_0/n 0.32fF
C274 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C275 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/k 0.21fF
C276 ffipg_0/pggen_0/xor_0/w_n3_4# x1in 0.06fF
C277 ffipg_2/k sumffo_2/xor_0/a_10_10# 0.12fF
C278 sumffo_0/xor_0/inv_0/w_0_6# ffipg_0/k 0.06fF
C279 cla_2/p0 ffipg_3/k 0.06fF
C280 gnd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C281 cla_0/g0 nand_2/b 0.13fF
C282 cla_2/p1 ffipg_3/pggen_0/nor_0/w_0_0# 0.05fF
C283 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C284 cla_0/l ffipg_2/k 0.10fF
C285 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C286 ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C287 ffipg_1/k y2in 0.07fF
C288 gnd sumffo_0/xor_0/w_n3_4# 0.12fF
C289 inv_8/w_0_6# inv_8/in 0.10fF
C290 cla_2/l inv_7/w_0_6# 0.06fF
C291 inv_0/op inv_0/in 0.04fF
C292 cla_0/l cla_0/n 0.25fF
C293 cin sumffo_3/xor_0/a_10_10# 0.04fF
C294 nor_1/w_0_0# inv_1/in 0.11fF
C295 gnd inv_4/op 0.58fF
C296 ffipg_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C297 inv_7/op gnd 0.27fF
C298 y4in gnd 1.76fF
C299 cla_2/nor_1/w_0_0# cla_2/inv_0/in 0.05fF
C300 ffipg_1/pggen_0/xor_0/a_10_10# y2in 0.12fF
C301 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C302 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C303 gnd inv_4/in 0.33fF
C304 inv_7/w_0_6# inv_7/in 0.10fF
C305 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C306 x3in cla_2/p0 0.22fF
C307 x4in ffipg_3/k 0.46fF
C308 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C309 cla_0/inv_0/op cla_0/nand_0/w_0_0# 0.06fF
C310 cla_0/l inv_7/w_0_6# 0.06fF
C311 inv_0/op cla_0/g0 0.32fF
C312 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C313 cla_1/n inv_4/in 0.02fF
C314 cla_2/inv_0/w_0_6# gnd 0.06fF
C315 cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# 0.04fF
C316 y4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C317 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C318 gnd sumffo_1/xor_0/inv_1/w_0_6# 0.06fF
C319 cla_2/p0 cla_2/p1 0.24fF
C320 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C321 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C322 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C323 ffipg_1/pggen_0/xor_0/inv_1/op y2in 0.22fF
C324 gnd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C325 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C326 sumffo_0/xor_0/op sumffo_0/xor_0/inv_1/op 0.52fF
C327 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C328 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C329 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C330 x1in ffipg_0/k 0.46fF
C331 gnd sumffo_0/xor_0/a_10_10# 0.93fF
C332 x2in ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C333 inv_8/w_0_6# cin 0.06fF
C334 inv_8/in gnd 0.43fF
C335 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.36fF
C336 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# x2in 0.06fF
C337 cla_0/l cla_0/nor_1/w_0_0# 0.02fF
C338 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C339 gnd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C340 x4in cla_2/p1 0.22fF
C341 ffipg_2/pggen_0/nand_0/w_0_0# cla_0/l 0.04fF
C342 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/op 0.06fF
C343 cla_0/inv_0/op nand_2/b 0.09fF
C344 ffipg_2/pggen_0/xor_0/inv_1/op y3in 0.22fF
C345 cla_0/nor_0/w_0_0# cla_0/l 0.05fF
C346 cla_0/n ffipg_2/k 0.06fF
C347 gnd ffipg_1/pggen_0/nand_0/a_13_n26# 0.01fF
C348 x1in ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C349 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C350 cla_1/inv_0/in cla_1/inv_0/op 0.04fF
C351 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C352 cla_2/g1 cla_2/p1 0.00fF
C353 cla_2/l inv_5/w_0_6# 0.08fF
C354 cin sumffo_0/xor_0/inv_0/op 0.20fF
C355 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C356 cla_2/l gnd 0.61fF
C357 gnd sumffo_1/xor_0/inv_1/op 0.35fF
C358 sumffo_3/xor_0/inv_1/w_0_6# ffipg_3/k 0.23fF
C359 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C360 cla_0/l cla_1/l 0.08fF
C361 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/op 0.02fF
C362 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C363 ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k 0.06fF
C364 gnd y1in 1.77fF
C365 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/a_10_10# 0.16fF
C366 gnd sumffo_2/xor_0/a_10_10# 0.93fF
C367 gnd inv_7/in 0.43fF
C368 sumffo_0/xor_0/op sumffo_0/xor_0/w_n3_4# 0.02fF
C369 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k 0.52fF
C370 nor_2/w_0_0# nor_2/b 0.06fF
C371 cla_0/inv_0/w_0_6# gnd 0.06fF
C372 sumffo_3/xor_0/inv_0/op ffipg_3/k 0.20fF
C373 x4in y4in 0.73fF
C374 inv_1/op ffipg_2/k 0.09fF
C375 cla_0/l gnd 3.30fF
C376 nor_0/a y1in 0.03fF
C377 cin gnd 1.53fF
C378 cla_0/l cla_1/nor_0/w_0_0# 0.01fF
C379 ffipg_2/pggen_0/xor_0/inv_0/op y3in 0.20fF
C380 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/k 0.45fF
C381 gnd sumffo_2/xor_0/w_n3_4# 0.12fF
C382 cla_2/g1 y4in 0.13fF
C383 cla_0/l nor_0/a 0.16fF
C384 ffipg_0/pggen_0/nor_0/w_0_0# y1in 0.06fF
C385 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C386 cla_1/n cla_0/l 0.13fF
C387 y4in ffipg_3/pggen_0/xor_0/inv_0/op 0.20fF
C388 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C389 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C390 inv_9/in gnd 0.33fF
C391 cla_1/p0 y2in 0.03fF
C392 inv_8/in nor_4/a 0.04fF
C393 nor_0/w_0_0# cinbar 0.06fF
C394 gnd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C395 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C396 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C397 ffipg_1/pggen_0/nand_0/w_0_0# y2in 0.06fF
C398 inv_3/in inv_3/w_0_6# 0.10fF
C399 cla_0/l inv_2/w_0_6# 0.06fF
C400 cin inv_0/in 0.07fF
C401 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# gnd 0.11fF
C402 cla_2/inv_0/in gnd 0.34fF
C403 cin inv_2/w_0_6# 0.06fF
C404 x4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C405 cla_0/g0 y1in 0.13fF
C406 cla_1/nand_0/a_13_n26# gnd 0.01fF
C407 cin ffipg_1/k 0.06fF
C408 ffipg_2/pggen_0/xor_0/a_10_10# y3in 0.12fF
C409 cla_2/l cla_2/p0 0.16fF
C410 sumffo_0/xor_0/op sumffo_0/xor_0/a_10_10# 0.45fF
C411 cla_2/nor_1/w_0_0# gnd 0.31fF
C412 cla_0/g0 cla_0/l 0.14fF
C413 gnd inv_3/in 0.47fF
C414 cla_0/g0 cin 0.08fF
C415 cin sumffo_1/xor_0/a_38_n43# 0.01fF
C416 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C417 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C418 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C419 cla_2/inv_0/op gnd 0.27fF
C420 cla_0/n inv_3/w_0_6# 0.16fF
C421 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k 0.52fF
C422 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C423 x3in ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C424 cla_1/l cla_0/n 0.07fF
C425 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C426 inv_2/in nor_1/b 0.04fF
C427 cla_0/l cla_2/p0 0.44fF
C428 gnd ffipg_2/k 0.64fF
C429 cla_0/n inv_5/w_0_6# 0.06fF
C430 gnd sumffo_3/xor_0/a_10_10# 0.93fF
C431 cin sumffo_3/xor_0/inv_1/op 0.04fF
C432 cla_0/n gnd 1.18fF
C433 gnd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C434 sumffo_3/xor_0/inv_0/op inv_4/op 0.27fF
C435 cla_2/l nor_3/b 0.10fF
C436 nand_2/b inv_2/in 0.34fF
C437 x1in y1in 0.73fF
C438 gnd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C439 cin sumffo_1/xor_0/a_10_10# 0.06fF
C440 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/op 0.06fF
C441 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C442 gnd sumffo_3/xor_0/w_n3_4# 0.12fF
C443 gnd inv_7/w_0_6# 0.15fF
C444 inv_9/in nor_4/a 0.02fF
C445 ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C446 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# gnd 0.09fF
C447 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C448 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_0/w_0_6# 0.03fF
C449 ffipg_0/pggen_0/xor_0/inv_0/op y1in 0.20fF
C450 x2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C451 gnd inv_1/op 0.58fF
C452 cla_0/l cla_2/g1 0.26fF
C453 nor_0/w_0_0# nand_2/b 0.04fF
C454 x3in ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C455 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.15fF
C456 cla_0/n nor_1/w_0_0# 0.06fF
C457 gnd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C458 inv_9/in nor_4/w_0_0# 0.11fF
C459 inv_4/op nor_2/w_0_0# 0.03fF
C460 x3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C461 inv_8/w_0_6# gnd 0.15fF
C462 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C463 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C464 cla_0/inv_0/op cla_0/l 0.35fF
C465 inv_4/in nor_2/w_0_0# 0.11fF
C466 x4in ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C467 ffipg_0/pggen_0/xor_0/inv_1/op y1in 0.22fF
C468 cla_0/nor_1/w_0_0# gnd 0.31fF
C469 cla_2/p0 ffipg_2/k 0.05fF
C470 ffipg_2/pggen_0/nand_0/w_0_0# gnd 0.10fF
C471 cla_0/nor_0/w_0_0# gnd 0.31fF
C472 ffipg_3/pggen_0/xor_0/inv_1/op y4in 0.22fF
C473 x3in y3in 0.73fF
C474 inv_9/in cout 0.04fF
C475 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C476 cla_2/nor_0/w_0_0# gnd 0.31fF
C477 nor_0/w_0_0# inv_0/op 0.10fF
C478 y4in ffipg_3/pggen_0/xor_0/a_10_10# 0.12fF
C479 cla_2/g1 cla_2/inv_0/in 0.04fF
C480 ffipg_0/pggen_0/xor_0/a_10_10# y1in 0.12fF
C481 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C482 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C483 inv_1/op nor_1/w_0_0# 0.03fF
C484 cla_1/l inv_3/w_0_6# 0.06fF
C485 gnd sumffo_0/xor_0/inv_0/op 0.36fF
C486 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C487 cla_0/l cla_1/inv_0/in 0.23fF
C488 ffipg_0/k cinbar 0.06fF
C489 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C490 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C491 gnd inv_3/w_0_6# 0.17fF
C492 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# 0.16fF
C493 cla_0/l cla_1/nand_0/w_0_0# 0.06fF
C494 y4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C495 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C496 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C497 cla_2/g1 cla_2/inv_0/op 0.35fF
C498 cla_1/l gnd 0.40fF
C499 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/op 0.06fF
C500 cla_0/l cla_1/p0 0.09fF
C501 x2in gnd 1.24fF
C502 gnd inv_5/w_0_6# 0.42fF
C503 cla_0/l ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C504 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C505 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C506 ffipg_1/pggen_0/nor_0/w_0_0# x2in 0.06fF
C507 ffipg_3/k ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C508 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/xor_0/inv_0/op 0.03fF
C509 ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C510 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C511 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/a_10_10# 0.16fF
C512 ffipg_1/pggen_0/nor_0/w_0_0# gnd 0.11fF
C513 gnd inv_6/in 0.33fF
C514 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C515 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C516 cla_1/nor_0/w_0_0# gnd 0.31fF
C517 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/k 0.02fF
C518 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C519 gnd nor_0/a 0.58fF
C520 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# x1in 0.06fF
C521 cla_1/n gnd 0.52fF
C522 inv_8/w_0_6# nor_4/a 0.03fF
C523 gnd ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C524 ffipg_2/pggen_0/nand_0/w_0_0# cla_2/p0 0.24fF
C525 ffipg_0/pggen_0/nor_0/w_0_0# gnd 0.11fF
C526 inv_9/in nor_4/b 0.16fF
C527 gnd inv_0/in 0.30fF
C528 sumffo_0/xor_0/inv_0/w_0_6# gnd 0.11fF
C529 x2in ffipg_1/k 0.46fF
C530 cla_2/nor_0/w_0_0# cla_2/p0 0.06fF
C531 gnd inv_2/w_0_6# 0.17fF
C532 gnd ffipg_1/k 0.76fF
C533 gnd nor_1/w_0_0# 0.17fF
C534 ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C535 ffipg_1/pggen_0/nor_0/w_0_0# ffipg_1/k 0.21fF
C536 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C537 inv_0/in nor_0/a 0.02fF
C538 gnd ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C539 gnd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C540 cla_0/g0 gnd 1.23fF
C541 ffipg_1/k nor_0/a 0.06fF
C542 cla_2/p1 ffipg_3/k 0.05fF
C543 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C544 inv_1/in nor_1/b 0.16fF
C545 inv_4/in nor_2/b 0.16fF
C546 cla_2/p0 cla_1/l 0.02fF
C547 cla_1/p0 ffipg_2/k 0.06fF
C548 cla_0/g0 nor_0/a 0.57fF
C549 cin sumffo_3/xor_0/a_38_n43# 0.01fF
C550 cla_1/inv_0/w_0_6# cla_1/inv_0/op 0.03fF
C551 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C552 cla_2/p0 gnd 1.12fF
C553 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C554 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C555 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C556 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C557 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C558 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C559 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C560 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C561 y4in Gnd 2.72fF
C562 x4in Gnd 2.80fF
C563 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C564 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C565 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C566 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C567 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C568 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C569 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C570 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C571 y3in Gnd 2.72fF
C572 x3in Gnd 2.80fF
C573 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C574 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C575 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C576 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C577 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C578 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C579 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C580 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C581 y2in Gnd 2.72fF
C582 x2in Gnd 2.80fF
C583 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C584 cout Gnd 0.19fF
C585 inv_9/in Gnd 0.23fF
C586 nor_4/w_0_0# Gnd 1.81fF
C587 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C588 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C589 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C590 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C591 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C592 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C593 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C594 y1in Gnd 2.72fF
C595 x1in Gnd 2.80fF
C596 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C597 nor_4/a Gnd 0.59fF
C598 inv_8/in Gnd 0.22fF
C599 inv_8/w_0_6# Gnd 1.40fF
C600 inv_7/in Gnd 0.22fF
C601 inv_7/w_0_6# Gnd 1.40fF
C602 nor_4/b Gnd 0.32fF
C603 nor_3/b Gnd 0.77fF
C604 inv_5/in Gnd 0.22fF
C605 inv_5/w_0_6# Gnd 1.40fF
C606 cla_2/n Gnd 0.36fF
C607 inv_6/in Gnd 0.23fF
C608 nor_3/w_0_0# Gnd 1.81fF
C609 cla_1/n Gnd 0.36fF
C610 inv_4/in Gnd 0.23fF
C611 nor_2/w_0_0# Gnd 1.81fF
C612 cla_0/n Gnd 1.34fF
C613 nor_2/b Gnd 0.82fF
C614 inv_3/in Gnd 0.22fF
C615 inv_3/w_0_6# Gnd 1.40fF
C616 cinbar Gnd 1.21fF
C617 nor_0/a Gnd 2.07fF
C618 nor_1/b Gnd 1.05fF
C619 inv_2/in Gnd 0.22fF
C620 inv_2/w_0_6# Gnd 1.40fF
C621 inv_1/in Gnd 0.23fF
C622 nor_1/w_0_0# Gnd 1.81fF
C623 inv_0/in Gnd 0.23fF
C624 sumffo_3/xor_0/op Gnd 0.06fF
C625 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C626 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C627 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C628 ffipg_3/k Gnd 2.89fF
C629 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C630 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C631 inv_4/op Gnd 1.37fF
C632 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C633 sumffo_1/xor_0/op Gnd 0.06fF
C634 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C635 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C636 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C637 nand_2/b Gnd 2.33fF
C638 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C639 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C640 ffipg_1/k Gnd 2.78fF
C641 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C642 sumffo_2/xor_0/op Gnd 0.06fF
C643 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C644 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C645 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C646 ffipg_2/k Gnd 2.89fF
C647 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C648 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C649 inv_1/op Gnd 1.30fF
C650 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C651 sumffo_0/xor_0/op Gnd 0.06fF
C652 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C653 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C654 gnd Gnd 32.08fF
C655 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C656 cin Gnd 7.80fF
C657 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C658 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C659 ffipg_0/k Gnd 1.49fF
C660 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C661 cla_2/p1 Gnd 1.09fF
C662 cla_2/nor_1/w_0_0# Gnd 1.23fF
C663 cla_2/nor_0/w_0_0# Gnd 1.23fF
C664 cla_2/inv_0/in Gnd 0.27fF
C665 cla_2/inv_0/w_0_6# Gnd 0.58fF
C666 cla_2/g1 Gnd 0.59fF
C667 cla_2/inv_0/op Gnd 0.26fF
C668 cla_2/nand_0/w_0_0# Gnd 0.82fF
C669 cla_2/p0 Gnd 0.38fF
C670 cla_1/nor_1/w_0_0# Gnd 1.23fF
C671 cla_1/l Gnd 0.30fF
C672 cla_1/nor_0/w_0_0# Gnd 1.23fF
C673 cla_1/inv_0/in Gnd 0.27fF
C674 cla_1/inv_0/w_0_6# Gnd 0.58fF
C675 cla_1/inv_0/op Gnd 0.26fF
C676 cla_1/nand_0/w_0_0# Gnd 0.82fF
C677 inv_7/op Gnd 0.26fF
C678 cla_1/p0 Gnd 2.28fF
C679 cla_0/nor_1/w_0_0# Gnd 1.23fF
C680 cla_0/l Gnd 3.41fF
C681 cla_0/nor_0/w_0_0# Gnd 1.23fF
C682 cla_0/inv_0/in Gnd 0.27fF
C683 cla_0/inv_0/w_0_6# Gnd 0.58fF
C684 cla_0/inv_0/op Gnd 0.26fF
C685 cla_0/nand_0/w_0_0# Gnd 0.82fF
C686 cla_2/l Gnd 0.25fF
C687 cla_0/g0 Gnd 1.40fF
C688 inv_0/op Gnd 0.23fF
C689 nor_0/w_0_0# Gnd 2.63fF
