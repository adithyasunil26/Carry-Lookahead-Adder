* SPICE3 file created from ffipgarrcla.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 vdd nand_5/a inv_1/in inv_1/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_1/in cla_0/l vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_1/in nand_5/a nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_2/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_0/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_2/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# nand_5/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd inv_7/op inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in nand_5/a vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in inv_7/op nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_0/g0 ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_0/g0 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1059 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1060 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1061 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1062 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1063 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1064 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 nor_0/a ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1069 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 gnd ffipgarr_0/ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1071 nor_0/a ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1073 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1074 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1076 ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1077 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1078 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 ffipgarr_0/ffipg_0/ffi_0/nand_1/a clk ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1081 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1082 ffipgarr_0/ffipg_0/ffi_0/nand_3/a y1in vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 ffipgarr_0/ffipg_0/ffi_0/nand_3/a clk ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1084 ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1086 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1088 ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1089 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1090 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1094 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1096 ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1097 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1098 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1101 vdd ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1102 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1107 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1108 ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1109 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1110 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1112 ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1113 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1114 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 ffipgarr_0/ffipg_0/ffi_1/nand_1/a clk ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1117 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1118 ffipgarr_0/ffipg_0/ffi_1/nand_3/a x1in vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 ffipgarr_0/ffipg_0/ffi_1/nand_3/a clk ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1122 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1124 ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1125 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1126 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1128 ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1129 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1130 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1133 vdd ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1134 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1136 ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1137 vdd ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1138 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1140 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1141 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1145 vdd ffipgarr_0/ffipg_1/ffi_0/q cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1146 cla_1/g0 ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1153 sumffo_1/k ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1154 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1155 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1156 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op sumffo_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 cla_1/p0 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1161 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 gnd ffipgarr_0/ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1163 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1165 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1166 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1168 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1169 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1170 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ffipgarr_0/ffipg_1/ffi_0/nand_1/a clk ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1172 ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1173 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1174 ffipgarr_0/ffipg_1/ffi_0/nand_3/a y2in vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 ffipgarr_0/ffipg_1/ffi_0/nand_3/a clk ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1176 ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1177 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1178 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1181 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1182 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1184 ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1185 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1186 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1188 ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1189 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1190 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1192 ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1193 vdd ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1194 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1201 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1202 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1204 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1205 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1206 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipgarr_0/ffipg_1/ffi_1/nand_1/a clk ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1208 ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1209 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1210 ffipgarr_0/ffipg_1/ffi_1/nand_3/a x2in vdd ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 ffipgarr_0/ffipg_1/ffi_1/nand_3/a clk ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1212 ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1213 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1214 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1216 ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1217 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1218 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1221 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1222 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1224 ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1225 vdd ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1226 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1228 ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1229 vdd ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1230 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1232 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1233 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1235 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1236 ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1237 vdd ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1238 cla_2/g0 ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 cla_2/g0 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1240 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1241 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1245 sumffo_2/k ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1246 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1247 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1248 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op sumffo_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1253 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 gnd ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1255 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1257 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1258 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1260 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1261 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1262 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 ffipgarr_0/ffipg_2/ffi_0/nand_1/a clk ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1264 ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1265 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1266 ffipgarr_0/ffipg_2/ffi_0/nand_3/a y3in vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 ffipgarr_0/ffipg_2/ffi_0/nand_3/a clk ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1268 ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1269 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1270 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1272 ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1273 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1274 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1276 ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1277 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1278 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1280 ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1281 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1282 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1284 ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1285 vdd ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1286 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1288 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1289 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1293 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1294 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1297 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1298 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 ffipgarr_0/ffipg_2/ffi_1/nand_1/a clk ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1301 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1302 ffipgarr_0/ffipg_2/ffi_1/nand_3/a x3in vdd ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 ffipgarr_0/ffipg_2/ffi_1/nand_3/a clk ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1304 ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1305 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1306 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1308 ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1309 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1310 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1313 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1314 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1316 ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1317 vdd ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1318 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1320 ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1321 vdd ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1322 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1325 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1326 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1327 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1328 ffipgarr_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1329 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1330 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/a vdd ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipgarr_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 vdd clk ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/inv_0/op vdd ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 ffipgarr_0/ffi_0/nand_1/a clk ffipgarr_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipgarr_0/ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1337 vdd clk ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1338 ffipgarr_0/ffi_0/nand_3/a cinin vdd ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 ffipgarr_0/ffi_0/nand_3/a clk ffipgarr_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 ffipgarr_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1341 vdd ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1342 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/a vdd ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1344 ffipgarr_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1345 vdd ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1346 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_3/b vdd ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1348 ffipgarr_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1349 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1350 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/inv_1/op vdd ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1352 ffipgarr_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 vdd nand_5/a nor_0/b ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 nor_0/b ffipgarr_0/ffi_0/nand_6/a vdd ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 nor_0/b nand_5/a ffipgarr_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipgarr_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 vdd nor_0/b nand_5/a ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 nand_5/a ffipgarr_0/ffi_0/nand_7/a vdd ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 nand_5/a nor_0/b ffipgarr_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipgarr_0/ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1361 ffipgarr_0/ffi_0/inv_0/op cinin vdd ffipgarr_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1362 ffipgarr_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1363 ffipgarr_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 vdd ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 cla_2/g1 ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1369 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1370 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1371 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1373 sumffo_3/k ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1374 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1375 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1376 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1381 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 gnd ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1383 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1385 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1386 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipgarr_0/ffipg_3/ffi_0/nand_1/a clk ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipgarr_0/ffipg_3/ffi_0/nand_3/a y4in vdd ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipgarr_0/ffipg_3/ffi_0/nand_3/a clk ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 vdd ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1417 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1418 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1419 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1421 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1422 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1425 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1426 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1427 ffipgarr_0/ffipg_3/ffi_1/nand_1/a clk ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1428 ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1429 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1430 ffipgarr_0/ffipg_3/ffi_1/nand_3/a x4in vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 ffipgarr_0/ffipg_3/ffi_1/nand_3/a clk ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1433 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1434 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1436 ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1437 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1438 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1440 ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1441 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1442 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1443 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1444 ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1445 vdd ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1446 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1448 ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1449 vdd ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1450 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1451 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1452 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1453 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1455 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1456 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1457 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1458 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1459 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1460 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1461 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1463 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1465 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1467 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1469 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1470 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a vdd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op vdd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1479 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1480 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 vdd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a vdd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 vdd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b vdd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 sumffo_0/ffo_0/nand_7/a clk vdd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 vdd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a vdd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 vdd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 z1o sumffo_0/ffo_0/nand_7/a vdd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1503 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1504 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1505 sumffo_0/ffo_0/nand_0/b clk vdd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 sumffo_0/xor_0/inv_0/op sumffo_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1507 sumffo_0/xor_0/inv_0/op sumffo_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1508 sumffo_0/xor_0/inv_1/op nand_5/a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1509 sumffo_0/xor_0/inv_1/op nand_5/a vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 vdd nand_5/a sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1511 sumffo_0/ffo_0/d nand_5/a sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1512 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1513 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1514 sumffo_0/xor_0/a_10_n43# sumffo_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1515 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 sumffo_0/xor_0/a_10_10# sumffo_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1520 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a vdd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1522 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1523 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1524 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op vdd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1527 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1528 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1529 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1530 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1531 vdd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1532 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a vdd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1534 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1535 vdd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1536 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b vdd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1538 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 sumffo_2/ffo_0/nand_7/a clk vdd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 vdd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a vdd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 vdd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 z3o sumffo_2/ffo_0/nand_7/a vdd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1551 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1552 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1553 sumffo_2/ffo_0/nand_0/b clk vdd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 sumffo_2/xor_0/inv_0/op sumffo_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1555 sumffo_2/xor_0/inv_0/op sumffo_2/k vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1556 sumffo_2/xor_0/inv_1/op inv_2/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1557 sumffo_2/xor_0/inv_1/op inv_2/op vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 vdd inv_2/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1559 sumffo_2/ffo_0/d inv_2/op sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1560 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1561 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1562 sumffo_2/xor_0/a_10_n43# sumffo_2/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 sumffo_2/xor_0/a_10_10# sumffo_2/k vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a vdd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1571 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1572 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op vdd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1573 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 vdd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a vdd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 vdd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b vdd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 sumffo_1/ffo_0/nand_7/a clk vdd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 vdd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a vdd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 vdd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 z2o sumffo_1/ffo_0/nand_7/a vdd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1599 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1600 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1601 sumffo_1/ffo_0/nand_0/b clk vdd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 sumffo_1/xor_0/inv_0/op sumffo_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1603 sumffo_1/xor_0/inv_0/op sumffo_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1604 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1605 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1607 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1608 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1609 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1610 sumffo_1/xor_0/a_10_n43# sumffo_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1611 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 sumffo_1/xor_0/a_10_10# sumffo_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1614 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a vdd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op vdd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 vdd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a vdd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 vdd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b vdd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 sumffo_3/ffo_0/nand_7/a clk vdd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 vdd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a vdd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1643 vdd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1644 z4o sumffo_3/ffo_0/nand_7/a vdd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1645 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1647 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1648 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1649 sumffo_3/ffo_0/nand_0/b clk vdd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 sumffo_3/xor_0/inv_0/op sumffo_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 sumffo_3/xor_0/inv_0/op sumffo_3/k vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 sumffo_3/xor_0/inv_1/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 sumffo_3/xor_0/inv_1/op inv_4/op vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 vdd inv_4/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 sumffo_3/ffo_0/d inv_4/op sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 sumffo_3/xor_0/a_10_n43# sumffo_3/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 sumffo_3/xor_0/a_10_10# sumffo_3/k vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1663 vdd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1664 ffo_0/nand_3/b ffo_0/nand_1/a vdd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1665 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1666 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 vdd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffo_0/nand_1/a ffo_0/inv_0/op vdd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 vdd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffo_0/nand_3/a ffo_0/d vdd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 vdd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffo_0/nand_1/b ffo_0/nand_3/a vdd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 vdd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffo_0/nand_6/a ffo_0/nand_3/b vdd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 vdd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffo_0/nand_7/a clk vdd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 vdd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffo_0/qbar ffo_0/nand_6/a vdd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 vdd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 couto ffo_0/nand_7/a vdd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1695 ffo_0/inv_0/op ffo_0/d vdd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1696 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1697 ffo_0/nand_0/b clk vdd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 nor_1/b inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 nor_1/b inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 inv_2/op inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1703 inv_2/op inv_2/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1704 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1705 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1706 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1707 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1708 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1709 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 inv_2/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1711 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 gnd nor_1/b inv_2/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1713 inv_2/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1714 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1715 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1716 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1717 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1719 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 nor_4/a inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1721 nor_4/a inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1723 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1724 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1725 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1726 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1727 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1728 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1729 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1730 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1731 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1732 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1733 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 nor_4/b inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 nor_4/b inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffo_0/d inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.34fF
C1 ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd 0.35fF
C2 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C3 ffo_0/nand_0/b ffo_0/d 0.40fF
C4 sumffo_3/k inv_4/op 0.09fF
C5 ffipgarr_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.06fF
C6 clk ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C7 sumffo_2/ffo_0/nand_0/w_0_0# cla_0/l 0.17fF
C8 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C9 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C10 nand_5/a clk 0.11fF
C11 gnd sumffo_1/ffo_0/inv_0/op 0.10fF
C12 cla_2/p0 cla_2/g0 0.16fF
C13 gnd ffo_0/nand_2/w_0_0# 0.00fF
C14 sumffo_3/ffo_0/nand_3/b vdd 0.39fF
C15 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C16 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.04fF
C17 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C18 vdd nor_0/w_0_0# 0.15fF
C19 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_1/a 0.04fF
C20 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C21 gnd ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.03fF
C22 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C23 gnd ffipgarr_0/ffi_0/nand_0/w_0_0# 0.00fF
C24 nor_0/b gnd 0.59fF
C25 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.06fF
C26 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C27 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_0/op 0.32fF
C28 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.03fF
C29 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C30 clk ffipgarr_0/ffi_0/nand_2/w_0_0# 0.06fF
C31 vdd sumffo_2/ffo_0/nand_0/w_0_0# 0.10fF
C32 vdd sumffo_0/ffo_0/nand_5/w_0_0# 0.10fF
C33 sumffo_3/ffo_0/inv_0/w_0_6# vdd 0.06fF
C34 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C35 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.15fF
C36 cla_0/n clk 0.12fF
C37 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# 0.06fF
C38 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C39 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# vdd 0.10fF
C40 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C41 vdd sumffo_1/ffo_0/nand_5/w_0_0# 0.10fF
C42 vdd sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C43 vdd sumffo_0/xor_0/a_10_10# 0.93fF
C44 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C45 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_3/b 0.00fF
C46 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/q 0.31fF
C47 gnd cla_0/g0 0.94fF
C48 sumffo_3/k cla_0/l 0.06fF
C49 cla_0/n sumffo_2/ffo_0/nand_3/a 0.07fF
C50 clk ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C51 inv_5/w_0_6# vdd 0.15fF
C52 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/inv_0/op 0.06fF
C53 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.04fF
C54 inv_8/w_0_6# inv_7/op 0.06fF
C55 gnd cla_1/p0 0.74fF
C56 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.13fF
C57 gnd ffo_0/nand_6/a 0.03fF
C58 vdd cla_1/nor_0/w_0_0# 0.32fF
C59 cla_0/n sumffo_2/ffo_0/nand_1/b 0.05fF
C60 cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C61 clk ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C62 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C63 gnd nor_1/b 0.10fF
C64 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C65 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a 0.13fF
C66 vdd sumffo_3/k 0.31fF
C67 vdd ffo_0/nand_4/w_0_0# 0.10fF
C68 clk ffo_0/nand_1/b 0.45fF
C69 inv_4/in nor_2/b 0.16fF
C70 gnd ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# 0.01fF
C71 ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd 0.22fF
C72 cla_1/nor_0/w_0_0# nand_2/b 0.01fF
C73 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# 0.04fF
C74 gnd ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.03fF
C75 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C76 sumffo_3/ffo_0/nand_6/a gnd 0.03fF
C77 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a 0.13fF
C78 vdd sumffo_0/sbar 0.28fF
C79 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.04fF
C80 vdd y4in 0.04fF
C81 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# clk 0.06fF
C82 gnd ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.03fF
C83 clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.13fF
C84 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.31fF
C85 clk ffo_0/nand_5/w_0_0# 0.06fF
C86 sumffo_3/xor_0/inv_0/op inv_4/op 0.20fF
C87 inv_2/op cla_0/l 0.06fF
C88 vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.17fF
C89 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.00fF
C90 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_0/op 0.06fF
C91 sumffo_0/xor_0/inv_1/w_0_6# sumffo_0/xor_0/inv_1/op 0.03fF
C92 gnd ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.26fF
C93 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C94 vdd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C95 vdd sumffo_2/k 0.29fF
C96 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.04fF
C97 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C98 clk nor_0/a 0.13fF
C99 ffo_0/nand_3/w_0_0# ffo_0/nand_3/b 0.06fF
C100 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.33fF
C101 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C102 x2in gnd 0.19fF
C103 inv_2/op vdd 0.34fF
C104 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# 0.04fF
C105 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C106 cla_1/inv_0/in cla_1/inv_0/op 0.04fF
C107 cla_0/nor_1/w_0_0# cla_0/g0 0.06fF
C108 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C109 gnd y2in 0.19fF
C110 vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.10fF
C111 ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd 0.30fF
C112 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C113 vdd sumffo_0/ffo_0/d 0.04fF
C114 gnd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.00fF
C115 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.10fF
C116 cla_1/p0 cla_0/nor_1/w_0_0# 0.06fF
C117 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C118 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/q 0.00fF
C119 sumffo_2/k nand_2/b 0.03fF
C120 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C121 clk ffo_0/inv_1/w_0_6# 0.06fF
C122 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C123 ffipgarr_0/ffipg_2/ffi_0/nand_1/b gnd 0.26fF
C124 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.04fF
C125 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C126 vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.34fF
C127 cla_0/n sumffo_2/ffo_0/nand_4/w_0_0# 0.24fF
C128 vdd x1in 0.04fF
C129 ffo_0/nand_3/w_0_0# vdd 0.11fF
C130 inv_2/op nand_2/b 0.10fF
C131 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/q 0.00fF
C132 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.15fF
C133 inv_3/in inv_3/w_0_6# 0.10fF
C134 gnd sumffo_0/ffo_0/nand_7/a 0.03fF
C135 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C136 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.04fF
C137 vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.10fF
C138 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# vdd 0.10fF
C139 vdd cla_2/p0 0.43fF
C140 nor_1/b nor_1/w_0_0# 0.06fF
C141 vdd ffipgarr_0/ffipg_3/ffi_0/qbar 0.33fF
C142 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C143 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C144 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.04fF
C145 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_0/op 0.06fF
C146 gnd cla_0/nand_0/w_0_0# 0.01fF
C147 vdd sumffo_3/xor_0/inv_0/op 0.15fF
C148 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op 1.63fF
C149 ffipgarr_0/ffi_0/nand_3/b gnd 0.35fF
C150 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.32fF
C151 nand_5/a ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.04fF
C152 vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C153 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.30fF
C154 cla_2/p0 nand_2/b 0.00fF
C155 z4o sumffo_3/ffo_0/nand_6/w_0_0# 0.06fF
C156 ffipgarr_0/ffi_0/nand_7/a nor_0/b 0.31fF
C157 ffo_0/nand_0/b vdd 0.15fF
C158 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.06fF
C159 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C160 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k 0.06fF
C161 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C162 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C163 gnd cla_2/nor_1/w_0_0# 0.01fF
C164 vdd sumffo_1/xor_0/inv_0/op 0.15fF
C165 cla_2/p1 cla_2/nor_0/w_0_0# 0.06fF
C166 cla_1/inv_0/w_0_6# cla_1/inv_0/op 0.03fF
C167 clk sumffo_3/ffo_0/nand_0/b 0.04fF
C168 nand_5/a inv_8/w_0_6# 0.57fF
C169 sumffo_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C170 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in 0.04fF
C171 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C172 cla_2/g0 cla_2/inv_0/in 0.16fF
C173 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.39fF
C174 vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C175 ffo_0/nand_7/a gnd 0.03fF
C176 vdd sumffo_3/sbar 0.28fF
C177 cla_0/n sumffo_2/ffo_0/nand_1/a 0.08fF
C178 nor_2/w_0_0# inv_4/op 0.03fF
C179 ffo_0/qbar ffo_0/nand_6/w_0_0# 0.04fF
C180 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C181 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C182 inv_3/w_0_6# nor_2/b 0.03fF
C183 vdd cla_2/n 0.28fF
C184 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C185 inv_5/w_0_6# inv_5/in 0.10fF
C186 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b 0.32fF
C187 x3in ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C188 vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C189 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.32fF
C190 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# vdd 0.93fF
C191 sumffo_1/xor_0/inv_0/op nand_2/b 0.20fF
C192 vdd sumffo_1/ffo_0/nand_3/w_0_0# 0.11fF
C193 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C194 cla_1/n gnd 0.08fF
C195 nor_0/b sumffo_0/k 0.09fF
C196 gnd cla_0/inv_0/in 0.35fF
C197 ffipgarr_0/ffipg_3/ffi_0/inv_1/op y4in 0.01fF
C198 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.13fF
C199 sumffo_1/ffo_0/inv_1/w_0_6# vdd 0.06fF
C200 vdd sumffo_2/xor_0/a_10_10# 0.93fF
C201 gnd ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.26fF
C202 ffipgarr_0/ffi_0/inv_0/w_0_6# cinin 0.06fF
C203 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_0/q 0.23fF
C204 clk sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C205 gnd sumffo_1/ffo_0/nand_3/a 0.03fF
C206 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/ffo_0/nand_7/a 0.06fF
C207 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C208 nand_5/a ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C209 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C210 cla_2/g1 cla_2/n 0.13fF
C211 cla_0/n cla_2/l 0.31fF
C212 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.04fF
C213 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.33fF
C214 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_1/op 0.52fF
C215 x4in ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C216 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.31fF
C217 x1in ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.01fF
C218 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.13fF
C219 sumffo_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C220 sumffo_1/ffo_0/nand_7/w_0_0# vdd 0.10fF
C221 gnd cinin 0.19fF
C222 ffo_0/nand_1/a gnd 0.03fF
C223 vdd ffipgarr_0/ffipg_2/ffi_1/q 1.35fF
C224 vdd ffo_0/d 0.19fF
C225 vdd sumffo_3/ffo_0/d 0.04fF
C226 nor_3/b cla_2/l 0.27fF
C227 sumffo_0/ffo_0/nand_6/a sumffo_0/sbar 0.00fF
C228 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# 0.04fF
C229 gnd ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.03fF
C230 sumffo_1/xor_0/inv_1/op gnd 0.20fF
C231 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C232 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.06fF
C233 sumffo_2/ffo_0/d gnd 0.37fF
C234 vdd sumffo_0/xor_0/inv_1/op 0.15fF
C235 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C236 inv_0/in vdd 0.09fF
C237 gnd sumffo_2/ffo_0/nand_7/a 0.03fF
C238 cla_2/g0 cla_0/l 0.08fF
C239 clk ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C240 nor_4/b inv_8/in 0.04fF
C241 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C242 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# vdd 0.10fF
C243 ffipgarr_0/ffipg_2/ffi_1/q nand_2/b 0.69fF
C244 gnd sumffo_2/ffo_0/inv_0/op 0.10fF
C245 nand_5/a nor_0/b 2.65fF
C246 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b 0.32fF
C247 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.06fF
C248 y2in ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C249 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.04fF
C250 gnd ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.15fF
C251 vdd nor_2/w_0_0# 0.15fF
C252 clk ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C253 vdd sumffo_0/xor_0/inv_1/w_0_6# 0.06fF
C254 inv_9/in ffo_0/d 0.04fF
C255 clk x4in 0.70fF
C256 gnd ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.22fF
C257 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.31fF
C258 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C259 ffo_0/nand_1/a ffo_0/nand_0/w_0_0# 0.04fF
C260 z4o gnd 0.52fF
C261 vdd sumffo_0/ffo_0/nand_2/w_0_0# 0.10fF
C262 vdd cla_2/g0 0.74fF
C263 gnd sumffo_2/ffo_0/nand_0/a_13_n26# 0.00fF
C264 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C265 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C266 inv_3/in gnd 0.36fF
C267 cla_0/nor_1/w_0_0# cla_0/inv_0/in 0.05fF
C268 nor_4/a vdd 0.15fF
C269 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_3/a 0.04fF
C270 ffipgarr_0/ffi_0/nand_6/w_0_0# nand_5/a 0.06fF
C271 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C272 nand_5/a cla_0/g0 0.05fF
C273 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# y4in 0.06fF
C274 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.15fF
C275 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a 0.00fF
C276 z4o sumffo_3/ffo_0/nand_7/a 0.00fF
C277 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.75fF
C278 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.04fF
C279 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C280 vdd y1in 0.04fF
C281 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C282 nand_5/a cla_1/p0 0.00fF
C283 vdd sumffo_1/ffo_0/nand_1/a 0.30fF
C284 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.03fF
C285 ffipgarr_0/ffi_0/inv_1/w_0_6# ffipgarr_0/ffi_0/inv_1/op 0.04fF
C286 gnd inv_1/w_0_6# 0.01fF
C287 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# sumffo_2/k 0.45fF
C288 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C289 clk sumffo_2/ffo_0/nand_1/b 0.45fF
C290 ffipgarr_0/ffi_0/nand_1/w_0_0# vdd 0.10fF
C291 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C292 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C293 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C294 cla_2/g1 cla_2/g0 0.44fF
C295 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.04fF
C296 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C297 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.06fF
C298 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_1/q 0.73fF
C299 sumffo_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C300 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.13fF
C301 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.04fF
C302 inv_9/in nor_4/a 0.02fF
C303 vdd z2o 0.28fF
C304 gnd ffo_0/inv_0/op 0.34fF
C305 sumffo_0/ffo_0/nand_7/w_0_0# z1o 0.04fF
C306 vdd cla_0/nor_0/w_0_0# 0.32fF
C307 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/inv_1/op 0.13fF
C308 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.04fF
C309 vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C310 vdd sumffo_2/ffo_0/nand_6/a 0.30fF
C311 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in 0.04fF
C312 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.04fF
C313 clk sumffo_1/ffo_0/d 0.05fF
C314 vdd ffipgarr_0/ffi_0/nand_7/w_0_0# 0.10fF
C315 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.06fF
C316 vdd ffipgarr_0/ffipg_0/ffi_1/q 1.35fF
C317 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C318 vdd cla_2/inv_0/in 0.05fF
C319 gnd ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.10fF
C320 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.06fF
C321 gnd ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.03fF
C322 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.31fF
C323 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C324 ffipgarr_0/ffipg_3/ffi_1/inv_0/op clk 0.32fF
C325 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.04fF
C326 inv_7/w_0_6# cla_0/l 0.06fF
C327 clk ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.07fF
C328 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C329 cla_0/n nor_1/b 0.37fF
C330 gnd nor_2/b 0.10fF
C331 inv_2/op inv_2/in 0.04fF
C332 ffo_0/inv_0/w_0_6# ffo_0/inv_0/op 0.03fF
C333 ffipgarr_0/ffipg_2/ffi_1/nand_1/b gnd 0.26fF
C334 sumffo_2/ffo_0/inv_0/w_0_6# sumffo_2/ffo_0/inv_0/op 0.03fF
C335 vdd inv_4/op 0.25fF
C336 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.04fF
C337 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C338 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk 0.07fF
C339 sumffo_2/k sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C340 gnd ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.03fF
C341 vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.10fF
C342 sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# 0.02fF
C343 vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.34fF
C344 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.00fF
C345 cla_2/g1 cla_2/inv_0/in 0.04fF
C346 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.30fF
C347 inv_7/w_0_6# vdd 0.20fF
C348 nor_0/b nor_0/a 0.39fF
C349 clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.13fF
C350 gnd ffipgarr_0/ffipg_0/ffi_0/qbar 0.34fF
C351 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C352 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q 0.27fF
C353 sumffo_0/xor_0/inv_0/w_0_6# sumffo_0/k 0.06fF
C354 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.06fF
C355 vdd ffipgarr_0/ffi_0/inv_0/op 0.17fF
C356 gnd ffipgarr_0/ffi_0/inv_1/op 0.22fF
C357 ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd 1.63fF
C358 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C359 cla_1/g0 cla_0/g0 0.18fF
C360 clk sumffo_1/ffo_0/nand_0/b 0.04fF
C361 clk sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C362 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.31fF
C363 gnd ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.10fF
C364 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.33fF
C365 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C366 cla_1/p0 cla_1/g0 1.76fF
C367 vdd sumffo_0/ffo_0/nand_3/a 0.30fF
C368 gnd ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.14fF
C369 vdd ffo_0/nand_3/b 0.39fF
C370 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/q 0.20fF
C371 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C372 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.31fF
C373 nor_0/a cla_0/g0 1.58fF
C374 gnd inv_8/in 0.13fF
C375 gnd ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# 0.01fF
C376 clk ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.32fF
C377 sumffo_1/xor_0/w_n3_4# vdd 0.12fF
C378 gnd ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.03fF
C379 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# y3in 0.06fF
C380 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.06fF
C381 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.00fF
C382 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.04fF
C383 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.10fF
C384 cla_1/p0 nor_0/a 0.24fF
C385 vdd cla_0/l 1.74fF
C386 couto vdd 0.28fF
C387 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.04fF
C388 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# 0.04fF
C389 vdd ffipgarr_0/ffipg_0/ffi_0/q 0.38fF
C390 inv_4/in nor_2/w_0_0# 0.11fF
C391 cla_1/n cla_1/nand_0/w_0_0# 0.04fF
C392 sumffo_3/ffo_0/nand_3/b gnd 0.35fF
C393 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/d 0.40fF
C394 x2in ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.06fF
C395 x1in ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C396 clk ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.32fF
C397 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# vdd 0.10fF
C398 vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.10fF
C399 nand_5/a ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.04fF
C400 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C401 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.04fF
C402 nand_2/b cla_0/l 0.46fF
C403 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.04fF
C404 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_0/op 0.32fF
C405 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# y4in 0.06fF
C406 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# vdd 0.10fF
C407 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.13fF
C408 ffipgarr_0/ffipg_0/ffi_0/q nand_2/b 0.90fF
C409 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.06fF
C410 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C411 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/d 0.40fF
C412 ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd 0.39fF
C413 sumffo_3/ffo_0/inv_0/w_0_6# gnd 0.01fF
C414 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.17fF
C415 cla_0/n cla_0/nand_0/w_0_0# 0.04fF
C416 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C417 sumffo_3/k ffipgarr_0/ffipg_3/ffi_0/q 0.07fF
C418 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C419 clk ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.06fF
C420 clk ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.32fF
C421 cla_2/nand_0/a_13_n26# gnd 0.01fF
C422 inv_1/in nor_1/b 0.04fF
C423 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.06fF
C424 vdd nand_2/b 0.82fF
C425 ffo_0/nand_6/a ffo_0/nand_6/w_0_0# 0.06fF
C426 cla_2/g1 vdd 0.35fF
C427 vdd ffipgarr_0/ffi_0/nand_3/w_0_0# 0.11fF
C428 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C429 inv_5/w_0_6# gnd 0.01fF
C430 inv_9/in vdd 0.09fF
C431 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C432 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/q 0.31fF
C433 vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.10fF
C434 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.06fF
C435 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.13fF
C436 sumffo_1/xor_0/inv_1/w_0_6# vdd 0.06fF
C437 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/b 0.31fF
C438 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C439 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C440 cla_1/p0 cla_1/l 0.16fF
C441 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C442 vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# 0.10fF
C443 clk sumffo_0/ffo_0/nand_0/b 0.04fF
C444 inv_7/in cla_2/l 0.13fF
C445 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.17fF
C446 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C447 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q 0.32fF
C448 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# 0.04fF
C449 sumffo_3/k gnd 0.35fF
C450 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/inv_1/op 0.45fF
C451 sumffo_0/ffo_0/nand_4/w_0_0# vdd 0.10fF
C452 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.10fF
C453 cla_2/p1 sumffo_3/k 0.05fF
C454 clk ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.06fF
C455 clk sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C456 sumffo_1/xor_0/inv_1/w_0_6# nand_2/b 0.23fF
C457 sumffo_2/xor_0/inv_1/op sumffo_2/k 0.06fF
C458 gnd sumffo_0/sbar 0.34fF
C459 gnd y4in 0.19fF
C460 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.06fF
C461 cla_0/n cla_1/n 0.09fF
C462 inv_4/in inv_4/op 0.04fF
C463 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/sbar 0.04fF
C464 cla_1/g0 cla_0/nand_0/w_0_0# 0.06fF
C465 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.11fF
C466 ffipgarr_0/ffi_0/nand_2/w_0_0# cinin 0.06fF
C467 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C468 gnd ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.10fF
C469 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/inv_0/op 0.06fF
C470 inv_2/op sumffo_2/xor_0/inv_1/op 0.22fF
C471 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.03fF
C472 ffo_0/nand_7/a ffo_0/nand_1/b 0.13fF
C473 gnd sumffo_2/k 0.35fF
C474 inv_7/op inv_8/in 0.13fF
C475 vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.10fF
C476 clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.13fF
C477 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.00fF
C478 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.13fF
C479 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op 0.06fF
C480 vdd sumffo_0/ffo_0/nand_1/b 0.31fF
C481 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.06fF
C482 ffo_0/nand_7/a ffo_0/nand_5/w_0_0# 0.04fF
C483 inv_2/op gnd 0.26fF
C484 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q 0.32fF
C485 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op 1.63fF
C486 vdd sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C487 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C488 ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd 0.15fF
C489 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.00fF
C490 gnd sumffo_0/ffo_0/d 0.37fF
C491 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op vdd 0.15fF
C492 sumffo_1/xor_0/w_n3_4# sumffo_1/k 0.06fF
C493 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.13fF
C494 sumffo_3/k ffipgarr_0/ffipg_3/ffi_1/q 0.46fF
C495 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# vdd 0.10fF
C496 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C497 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.00fF
C498 vdd nand_0/w_0_0# 0.10fF
C499 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C500 clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.13fF
C501 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C502 clk ffipgarr_0/ffi_0/nand_0/w_0_0# 0.06fF
C503 gnd ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.03fF
C504 gnd x1in 0.19fF
C505 vdd cla_1/nor_0/a_13_6# 0.01fF
C506 nor_3/w_0_0# cla_2/n 0.06fF
C507 vdd sumffo_1/ffo_0/inv_0/w_0_6# 0.08fF
C508 sumffo_1/ffo_0/nand_4/w_0_0# vdd 0.10fF
C509 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/qbar 0.00fF
C510 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C511 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.20fF
C512 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.04fF
C513 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C514 clk ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C515 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C516 cla_1/g0 cla_0/inv_0/in 0.04fF
C517 nand_5/a inv_1/w_0_6# 0.06fF
C518 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C519 sumffo_2/sbar z3o 0.32fF
C520 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.00fF
C521 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C522 vdd sumffo_1/k 0.26fF
C523 gnd cla_2/p0 0.74fF
C524 gnd ffipgarr_0/ffipg_3/ffi_0/qbar 0.34fF
C525 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 1.63fF
C526 vdd cla_0/inv_0/op 0.17fF
C527 sumffo_3/ffo_0/nand_0/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C528 cla_2/p1 cla_2/p0 0.24fF
C529 y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.04fF
C530 nand_2/b nand_0/w_0_0# 0.04fF
C531 inv_3/in cla_0/n 0.02fF
C532 inv_4/in vdd 0.09fF
C533 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# cla_2/g1 0.04fF
C534 nor_4/b nor_4/a 0.35fF
C535 clk cla_0/g0 0.10fF
C536 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C537 gnd ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.22fF
C538 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C539 cla_1/nor_0/a_13_6# nand_2/b 0.01fF
C540 sumffo_0/xor_0/w_n3_4# sumffo_0/k 0.06fF
C541 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C542 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.13fF
C543 vdd cla_0/nor_0/a_13_6# 0.01fF
C544 inv_5/in vdd 0.30fF
C545 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C546 clk ffo_0/nand_6/a 0.13fF
C547 ffo_0/nand_3/a ffo_0/nand_2/w_0_0# 0.04fF
C548 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d 0.04fF
C549 gnd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.00fF
C550 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.04fF
C551 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.33fF
C552 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_0/q 0.12fF
C553 vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.10fF
C554 gnd ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.14fF
C555 sumffo_1/k nand_2/b 0.51fF
C556 ffo_0/nand_0/b gnd 0.43fF
C557 vdd sumffo_0/ffo_0/nand_6/a 0.30fF
C558 x3in vdd 0.04fF
C559 vdd ffipgarr_0/ffi_0/nand_3/a 0.30fF
C560 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C561 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C562 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.00fF
C563 inv_0/op cla_0/g0 0.32fF
C564 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/w_0_0# 0.06fF
C565 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C566 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C567 z1o sumffo_0/ffo_0/nand_7/a 0.00fF
C568 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.04fF
C569 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.35fF
C570 gnd sumffo_3/sbar 0.34fF
C571 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.06fF
C572 cla_1/nand_0/a_13_n26# cla_0/l 0.01fF
C573 ffipgarr_0/ffi_0/nand_4/w_0_0# vdd 0.10fF
C574 clk ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.07fF
C575 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_0/qbar 0.06fF
C576 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C577 clk sumffo_3/ffo_0/nand_6/a 0.13fF
C578 gnd cla_2/n 0.22fF
C579 clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.13fF
C580 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.04fF
C581 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.04fF
C582 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/op 0.04fF
C583 inv_2/op nor_1/w_0_0# 0.03fF
C584 ffipgarr_0/ffi_0/nand_0/a_13_n26# gnd 0.01fF
C585 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.06fF
C586 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.06fF
C587 sumffo_3/ffo_0/nand_7/a sumffo_3/sbar 0.31fF
C588 vdd sumffo_3/ffo_0/nand_1/b 0.31fF
C589 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C590 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_1/w_0_6# 0.03fF
C591 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C592 ffo_0/qbar ffo_0/nand_6/a 0.00fF
C593 nand_5/a sumffo_0/xor_0/w_n3_4# 0.06fF
C594 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C595 cla_0/n nor_2/b 0.22fF
C596 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_1/b 0.04fF
C597 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# vdd 0.93fF
C598 ffo_0/nand_0/b ffo_0/nand_0/w_0_0# 0.06fF
C599 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.06fF
C600 vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C601 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/b 0.32fF
C602 vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C603 vdd y3in 0.04fF
C604 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C605 clk x2in 0.70fF
C606 nor_3/w_0_0# nor_4/a 0.03fF
C607 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C608 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C609 nand_5/a inv_8/in 0.00fF
C610 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C611 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C612 clk y2in 0.70fF
C613 vdd sumffo_2/ffo_0/nand_3/b 0.39fF
C614 ffipgarr_0/ffipg_2/ffi_1/q gnd 0.93fF
C615 gnd ffo_0/d 0.26fF
C616 gnd sumffo_3/ffo_0/d 0.37fF
C617 clk ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.06fF
C618 z3o sumffo_2/ffo_0/nand_6/w_0_0# 0.06fF
C619 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.45fF
C620 vdd inv_2/in 0.09fF
C621 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# 0.04fF
C622 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# vdd 0.10fF
C623 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C624 ffipgarr_0/ffipg_2/ffi_1/qbar vdd 0.33fF
C625 inv_3/w_0_6# cla_0/l 0.17fF
C626 inv_0/in gnd 0.24fF
C627 vdd sumffo_1/xor_0/a_10_10# 0.93fF
C628 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.75fF
C629 ffo_0/inv_0/w_0_6# ffo_0/d 0.06fF
C630 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.06fF
C631 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C632 vdd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C633 vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.34fF
C634 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C635 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C636 gnd ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# 0.01fF
C637 cla_2/g0 cla_1/nor_1/w_0_0# 0.02fF
C638 vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C639 inv_3/w_0_6# vdd 0.15fF
C640 inv_1/in inv_1/w_0_6# 0.10fF
C641 nand_5/a ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.04fF
C642 vdd sumffo_1/ffo_0/nand_2/w_0_0# 0.10fF
C643 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C644 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.31fF
C645 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.31fF
C646 gnd cla_2/g0 0.32fF
C647 sumffo_1/xor_0/a_10_10# nand_2/b 0.12fF
C648 vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.17fF
C649 cla_2/p1 cla_2/g0 0.35fF
C650 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.45fF
C651 nor_4/a gnd 0.15fF
C652 nor_4/b vdd 0.41fF
C653 nand_5/a sumffo_0/xor_0/a_10_10# 0.12fF
C654 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.17fF
C655 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.31fF
C656 inv_2/op sumffo_2/xor_0/inv_1/w_0_6# 0.23fF
C657 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C658 vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.34fF
C659 gnd y1in 0.19fF
C660 vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C661 gnd sumffo_1/ffo_0/nand_1/a 0.27fF
C662 cla_0/n sumffo_2/ffo_0/nand_0/w_0_0# 0.04fF
C663 sumffo_3/ffo_0/nand_1/a vdd 0.30fF
C664 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_1/b 0.31fF
C665 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.32fF
C666 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C667 inv_3/w_0_6# nand_2/b 0.06fF
C668 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_1/b 0.04fF
C669 ffipgarr_0/ffi_0/nand_1/a vdd 0.30fF
C670 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.30fF
C671 cla_2/p0 cla_1/inv_0/in 0.02fF
C672 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C673 vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C674 sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# 0.04fF
C675 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.04fF
C676 vdd sumffo_3/ffo_0/nand_6/w_0_0# 0.10fF
C677 gnd z2o 0.52fF
C678 vdd ffipgarr_0/ffipg_1/ffi_1/q 1.33fF
C679 inv_9/in nor_4/b 0.16fF
C680 sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# 0.04fF
C681 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/q 0.00fF
C682 inv_5/w_0_6# cla_0/n 0.06fF
C683 gnd sumffo_2/ffo_0/nand_6/a 0.03fF
C684 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C685 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# vdd 0.10fF
C686 vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.34fF
C687 gnd ffipgarr_0/ffipg_0/ffi_1/q 0.94fF
C688 gnd cla_2/inv_0/in 0.35fF
C689 ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd 0.30fF
C690 inv_5/w_0_6# nor_3/b 0.03fF
C691 cla_2/p1 cla_2/inv_0/in 0.02fF
C692 vdd ffipgarr_0/ffipg_2/ffi_0/qbar 0.33fF
C693 vdd ffipgarr_0/ffipg_1/ffi_0/q 0.38fF
C694 z4o sumffo_3/ffo_0/nand_7/w_0_0# 0.04fF
C695 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.06fF
C696 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.00fF
C697 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.06fF
C698 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.06fF
C699 cla_0/n sumffo_3/k 0.05fF
C700 ffo_0/nand_7/a ffo_0/qbar 0.31fF
C701 vdd sumffo_0/ffo_0/nand_3/w_0_0# 0.11fF
C702 gnd inv_4/op 0.21fF
C703 ffipgarr_0/ffi_0/inv_1/w_0_6# vdd 0.06fF
C704 clk cinin 0.70fF
C705 z2o sumffo_1/ffo_0/nand_6/a 0.31fF
C706 vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.10fF
C707 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C708 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C709 gnd ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.03fF
C710 ffipgarr_0/ffi_0/inv_0/w_0_6# ffipgarr_0/ffi_0/inv_0/op 0.03fF
C711 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C712 vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.10fF
C713 nor_0/w_0_0# nor_0/a 0.06fF
C714 vdd sumffo_3/ffo_0/nand_3/w_0_0# 0.11fF
C715 clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.13fF
C716 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_3/b 0.00fF
C717 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# vdd 0.10fF
C718 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.04fF
C719 gnd ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.14fF
C720 nor_3/w_0_0# vdd 0.17fF
C721 vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C722 nand_2/b ffipgarr_0/ffipg_1/ffi_0/q 0.32fF
C723 vdd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C724 sumffo_2/k sumffo_2/xor_0/inv_0/op 0.27fF
C725 gnd ffipgarr_0/ffi_0/inv_0/op 0.10fF
C726 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C727 vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.10fF
C728 ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd 0.22fF
C729 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.06fF
C730 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C731 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.06fF
C732 vdd ffipgarr_0/ffi_0/nand_6/a 0.30fF
C733 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/qbar 0.31fF
C734 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.39fF
C735 clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.13fF
C736 inv_2/op sumffo_2/xor_0/inv_0/op 0.20fF
C737 gnd sumffo_0/ffo_0/nand_3/a 0.03fF
C738 gnd ffo_0/nand_3/b 0.35fF
C739 vdd ffipgarr_0/ffipg_3/ffi_0/q 0.38fF
C740 clk ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.07fF
C741 cla_0/n inv_2/op 0.70fF
C742 vdd sumffo_2/ffo_0/nand_7/w_0_0# 0.10fF
C743 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b 0.13fF
C744 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/inv_0/op 0.03fF
C745 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.06fF
C746 vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.10fF
C747 gnd cla_0/l 0.88fF
C748 couto gnd 0.52fF
C749 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# 0.04fF
C750 vdd sumffo_2/xor_0/inv_1/op 0.15fF
C751 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.06fF
C752 gnd ffipgarr_0/ffipg_0/ffi_0/q 2.63fF
C753 vdd cla_2/nand_0/w_0_0# 0.10fF
C754 clk sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C755 vdd ffipgarr_0/ffi_0/inv_0/w_0_6# 0.06fF
C756 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C757 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.06fF
C758 sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d 0.52fF
C759 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C760 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a 0.31fF
C761 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C762 vdd cla_1/nor_1/w_0_0# 0.31fF
C763 x4in ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C764 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q 0.13fF
C765 ffipgarr_0/ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C766 vdd gnd 7.08fF
C767 vdd sumffo_1/ffo_0/nand_1/b 0.31fF
C768 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.45fF
C769 clk ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C770 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C771 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.31fF
C772 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C773 cla_2/p1 vdd 0.31fF
C774 ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd 0.35fF
C775 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C776 sumffo_2/k cla_1/g0 0.56fF
C777 vdd sumffo_3/ffo_0/nand_7/a 0.30fF
C778 cla_2/g1 cla_2/nand_0/w_0_0# 0.06fF
C779 cla_1/inv_0/in cla_2/g0 0.04fF
C780 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C781 ffo_0/inv_0/w_0_6# vdd 0.06fF
C782 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C783 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_1/b 0.04fF
C784 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.04fF
C785 vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C786 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.31fF
C787 clk ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.32fF
C788 gnd nand_2/b 1.54fF
C789 sumffo_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C790 ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd 0.39fF
C791 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C792 cla_2/g1 gnd 0.27fF
C793 inv_9/in gnd 0.24fF
C794 vdd sumffo_1/ffo_0/nand_6/a 0.30fF
C795 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.04fF
C796 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.13fF
C797 sumffo_1/k ffipgarr_0/ffipg_1/ffi_1/q 0.46fF
C798 cla_1/p0 cla_0/g0 0.33fF
C799 sumffo_2/ffo_0/nand_1/w_0_0# vdd 0.10fF
C800 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C801 sumffo_1/sbar sumffo_1/ffo_0/nand_7/w_0_0# 0.06fF
C802 cla_2/p1 cla_2/g1 0.17fF
C803 clk ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C804 vdd ffo_0/nand_0/w_0_0# 0.10fF
C805 sumffo_3/xor_0/a_10_10# sumffo_3/ffo_0/d 0.45fF
C806 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# vdd 0.10fF
C807 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C808 sumffo_2/ffo_0/nand_7/a z3o 0.00fF
C809 clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.13fF
C810 sumffo_1/k ffipgarr_0/ffipg_1/ffi_0/q 0.07fF
C811 cla_1/nand_0/w_0_0# cla_2/g0 0.06fF
C812 inv_7/w_0_6# inv_7/op 0.03fF
C813 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.32fF
C814 vdd ffipgarr_0/ffipg_3/ffi_1/q 1.35fF
C815 vdd sumffo_3/ffo_0/nand_1/w_0_0# 0.10fF
C816 cla_2/nor_0/w_0_0# cla_2/l 0.05fF
C817 cla_1/g0 cla_2/p0 0.32fF
C818 vdd sumffo_1/ffo_0/nand_3/b 0.39fF
C819 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/qbar 0.00fF
C820 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C821 sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d 0.06fF
C822 clk ffipgarr_0/ffi_0/inv_1/op 0.10fF
C823 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C824 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C825 nor_3/b cla_2/n 0.37fF
C826 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/b 0.31fF
C827 vdd cla_0/nor_1/w_0_0# 0.31fF
C828 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/q 0.20fF
C829 nand_5/a sumffo_0/xor_0/inv_1/op 0.22fF
C830 vdd sumffo_0/ffo_0/inv_0/op 0.17fF
C831 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# sumffo_2/k 0.01fF
C832 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C833 clk ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.32fF
C834 clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.13fF
C835 vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.10fF
C836 vdd nor_1/w_0_0# 0.15fF
C837 vdd sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C838 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_3/b 0.31fF
C839 ffo_0/nand_7/w_0_0# ffo_0/qbar 0.06fF
C840 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.30fF
C841 cla_2/inv_0/op cla_2/inv_0/in 0.04fF
C842 nand_5/a sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C843 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.15fF
C844 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C845 gnd sumffo_0/ffo_0/nand_1/b 0.26fF
C846 vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.10fF
C847 cla_0/nor_1/w_0_0# nand_2/b 0.02fF
C848 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.45fF
C849 gnd ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.22fF
C850 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C851 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.04fF
C852 clk ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C853 ffipgarr_0/ffi_0/nand_1/b vdd 0.31fF
C854 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.39fF
C855 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op gnd 0.17fF
C856 sumffo_0/k ffipgarr_0/ffipg_0/ffi_1/q 1.58fF
C857 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C858 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C859 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.31fF
C860 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.06fF
C861 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C862 z1o sumffo_0/sbar 0.32fF
C863 vdd inv_7/op 0.15fF
C864 vdd sumffo_0/ffo_0/nand_3/b 0.39fF
C865 cla_2/p1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C866 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C867 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.13fF
C868 sumffo_1/sbar z2o 0.32fF
C869 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.31fF
C870 clk sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C871 ffo_0/nand_0/b ffo_0/inv_1/w_0_6# 0.03fF
C872 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.04fF
C873 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# 0.04fF
C874 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C875 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.04fF
C876 gnd sumffo_1/k 0.35fF
C877 nor_0/w_0_0# inv_0/op 0.03fF
C878 gnd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.22fF
C879 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/w_0_0# 0.04fF
C880 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.11fF
C881 gnd cla_0/inv_0/op 0.15fF
C882 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# 0.04fF
C883 clk ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C884 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C885 inv_4/in gnd 0.24fF
C886 cla_2/p0 cla_1/l 0.02fF
C887 clk sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C888 clk sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C889 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C890 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C891 vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.10fF
C892 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.04fF
C893 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.45fF
C894 nand_5/a cla_0/nor_0/w_0_0# 0.01fF
C895 vdd ffipgarr_0/ffipg_3/ffi_1/qbar 0.33fF
C896 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/q 0.00fF
C897 ffipgarr_0/ffipg_2/ffi_1/q cla_1/g0 0.93fF
C898 inv_5/in gnd 0.17fF
C899 vdd sumffo_2/ffo_0/nand_5/w_0_0# 0.10fF
C900 nand_5/a ffipgarr_0/ffipg_0/ffi_1/q 0.02fF
C901 inv_4/op sumffo_3/xor_0/a_10_10# 0.12fF
C902 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_6/a 0.04fF
C903 gnd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.00fF
C904 nand_5/a ffipgarr_0/ffi_0/nand_7/w_0_0# 0.04fF
C905 ffipgarr_0/ffi_0/nand_7/a vdd 0.30fF
C906 gnd sumffo_0/ffo_0/nand_6/a 0.03fF
C907 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C908 vdd cla_1/inv_0/in 0.05fF
C909 x3in gnd 0.19fF
C910 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C911 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.06fF
C912 gnd ffipgarr_0/ffi_0/nand_3/a 0.03fF
C913 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.04fF
C914 sumffo_2/ffo_0/nand_0/b vdd 0.15fF
C915 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q 0.27fF
C916 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/qbar 0.00fF
C917 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C918 clk ffo_0/nand_4/w_0_0# 0.06fF
C919 vdd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C920 cla_1/nand_0/w_0_0# cla_0/l 0.08fF
C921 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/inv_1/w_0_6# 0.03fF
C922 sumffo_0/ffo_0/inv_0/w_0_6# sumffo_0/ffo_0/inv_0/op 0.03fF
C923 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C924 vdd sumffo_2/xor_0/inv_1/w_0_6# 0.06fF
C925 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C926 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C927 inv_0/in nor_0/a 0.02fF
C928 vdd cla_2/inv_0/op 0.17fF
C929 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.06fF
C930 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q 0.07fF
C931 clk y4in 0.64fF
C932 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d 0.04fF
C933 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.45fF
C934 sumffo_1/ffo_0/nand_4/w_0_0# sumffo_1/ffo_0/nand_3/b 0.06fF
C935 nor_4/w_0_0# ffo_0/d 0.03fF
C936 gnd sumffo_3/ffo_0/nand_1/b 0.26fF
C937 cla_1/g0 cla_2/g0 0.13fF
C938 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_1/op 0.08fF
C939 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# 0.04fF
C940 clk ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.32fF
C941 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.06fF
C942 cla_0/g0 cla_0/inv_0/in 0.16fF
C943 vdd cla_1/nand_0/w_0_0# 0.10fF
C944 vdd sumffo_0/k 0.31fF
C945 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C946 cla_1/p0 cla_0/inv_0/in 0.02fF
C947 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C948 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.31fF
C949 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# gnd 0.01fF
C950 gnd y3in 0.19fF
C951 cla_2/g1 cla_2/inv_0/op 0.35fF
C952 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b 0.32fF
C953 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.32fF
C954 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# vdd 0.06fF
C955 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.30fF
C956 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.04fF
C957 clk inv_2/op 1.02fF
C958 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# vdd 0.10fF
C959 vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.10fF
C960 gnd sumffo_2/ffo_0/nand_3/b 0.52fF
C961 clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.13fF
C962 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_1/q 0.73fF
C963 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.45fF
C964 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.06fF
C965 clk sumffo_0/ffo_0/d 0.25fF
C966 sumffo_1/sbar vdd 0.28fF
C967 vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.34fF
C968 nand_5/a cla_0/l 0.36fF
C969 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C970 vdd cla_1/inv_0/w_0_6# 0.06fF
C971 gnd inv_2/in 0.24fF
C972 vdd sumffo_3/xor_0/a_10_10# 0.93fF
C973 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.04fF
C974 nand_5/a ffipgarr_0/ffipg_0/ffi_0/q 0.02fF
C975 inv_6/in cla_2/n 0.02fF
C976 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.06fF
C977 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.00fF
C978 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.04fF
C979 clk x1in 0.70fF
C980 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.31fF
C981 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C982 ffipgarr_0/ffipg_2/ffi_1/qbar gnd 0.34fF
C983 nor_4/w_0_0# nor_4/a 0.06fF
C984 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C985 vdd sumffo_0/ffo_0/nand_6/w_0_0# 0.10fF
C986 vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.10fF
C987 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.04fF
C988 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/d 0.40fF
C989 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C990 nand_5/a vdd 1.48fF
C991 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.04fF
C992 nor_0/a cla_0/nor_0/w_0_0# 0.06fF
C993 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C994 ffipgarr_0/ffipg_3/ffi_1/inv_1/op x4in 0.01fF
C995 gnd ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.03fF
C996 cla_0/n cla_0/l 0.83fF
C997 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_3/b 0.04fF
C998 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.10fF
C999 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.04fF
C1000 nor_0/a ffipgarr_0/ffipg_0/ffi_1/q 0.22fF
C1001 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.07fF
C1002 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar 0.32fF
C1003 inv_3/w_0_6# gnd 0.01fF
C1004 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.39fF
C1005 inv_8/w_0_6# inv_8/in 0.10fF
C1006 ffipgarr_0/ffi_0/nand_2/w_0_0# vdd 0.10fF
C1007 gnd ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.10fF
C1008 sumffo_2/xor_0/w_n3_4# sumffo_2/k 0.06fF
C1009 vdd sumffo_2/xor_0/inv_0/op 0.15fF
C1010 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.32fF
C1011 clk ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C1012 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1013 ffipgarr_0/ffipg_2/ffi_0/q sumffo_2/k 0.07fF
C1014 clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.13fF
C1015 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.04fF
C1016 nor_4/b gnd 0.67fF
C1017 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C1018 gnd ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.26fF
C1019 clk ffo_0/nand_0/b 0.04fF
C1020 cla_0/n vdd 0.68fF
C1021 gnd ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.03fF
C1022 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# 0.04fF
C1023 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# cla_1/p0 0.05fF
C1024 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C1025 ffo_0/nand_1/b ffo_0/nand_3/b 0.32fF
C1026 sumffo_3/ffo_0/nand_1/a gnd 0.03fF
C1027 inv_2/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1028 ffo_0/nand_3/w_0_0# ffo_0/nand_3/a 0.06fF
C1029 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.04fF
C1030 ffipgarr_0/ffi_0/nand_1/a gnd 0.14fF
C1031 gnd ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.03fF
C1032 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.06fF
C1033 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1034 nor_3/b vdd 0.35fF
C1035 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C1036 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.04fF
C1037 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C1038 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.06fF
C1039 ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd 0.34fF
C1040 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/sbar 0.06fF
C1041 cla_0/n nand_2/b 0.05fF
C1042 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# vdd 0.10fF
C1043 nor_1/b inv_1/w_0_6# 0.03fF
C1044 gnd ffipgarr_0/ffipg_1/ffi_1/q 0.93fF
C1045 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1046 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.31fF
C1047 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.06fF
C1048 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.04fF
C1049 inv_2/in nor_1/w_0_0# 0.11fF
C1050 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C1051 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# gnd 0.00fF
C1052 gnd ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.03fF
C1053 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C1054 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.04fF
C1055 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C1056 vdd ffo_0/nand_1/b 0.31fF
C1057 ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd 0.03fF
C1058 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C1059 ffipgarr_0/ffipg_2/ffi_0/q cla_2/p0 0.03fF
C1060 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.04fF
C1061 nor_4/a inv_6/in 0.04fF
C1062 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C1063 vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C1064 sumffo_2/ffo_0/nand_2/w_0_0# cla_0/l 0.17fF
C1065 ffo_0/nand_3/a ffo_0/nand_0/b 0.13fF
C1066 gnd ffipgarr_0/ffipg_2/ffi_0/qbar 0.34fF
C1067 gnd ffipgarr_0/ffipg_1/ffi_0/q 2.58fF
C1068 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.04fF
C1069 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# vdd 0.06fF
C1070 nor_0/a cla_0/l 0.16fF
C1071 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C1072 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C1073 ffipgarr_0/ffipg_1/ffi_0/inv_1/op y2in 0.01fF
C1074 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.30fF
C1075 vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.10fF
C1076 cla_0/nand_0/a_13_n26# nand_2/b 0.00fF
C1077 vdd ffo_0/nand_5/w_0_0# 0.10fF
C1078 sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d 0.06fF
C1079 ffipgarr_0/ffipg_0/ffi_0/q nor_0/a 0.14fF
C1080 vdd cla_1/g0 0.49fF
C1081 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1082 clk sumffo_3/ffo_0/d 0.26fF
C1083 gnd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.00fF
C1084 inv_5/w_0_6# cla_2/l 0.29fF
C1085 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C1086 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C1087 vdd sumffo_2/ffo_0/nand_2/w_0_0# 0.10fF
C1088 y4in ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.04fF
C1089 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.04fF
C1090 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.04fF
C1091 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in 0.04fF
C1092 vdd nor_0/a 0.29fF
C1093 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.08fF
C1094 vdd ffipgarr_0/ffipg_0/ffi_1/qbar 0.33fF
C1095 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# x2in 0.06fF
C1096 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1097 inv_1/in cla_0/l 0.08fF
C1098 cla_1/g0 nand_2/b 1.65fF
C1099 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C1100 gnd ffipgarr_0/ffi_0/nand_6/a 0.03fF
C1101 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.33fF
C1102 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C1103 sumffo_0/ffo_0/nand_1/a vdd 0.30fF
C1104 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# sumffo_3/k 0.21fF
C1105 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.06fF
C1106 gnd ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.35fF
C1107 vdd sumffo_0/xor_0/inv_0/op 0.15fF
C1108 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_0/q 0.23fF
C1109 vdd sumffo_3/ffo_0/inv_0/op 0.17fF
C1110 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C1111 nor_0/b nor_0/w_0_0# 0.06fF
C1112 vdd ffo_0/inv_1/w_0_6# 0.06fF
C1113 nor_4/w_0_0# vdd 0.15fF
C1114 gnd ffipgarr_0/ffipg_3/ffi_0/q 2.62fF
C1115 nand_2/b nor_0/a 1.53fF
C1116 z2o sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C1117 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C1118 couto ffo_0/nand_6/w_0_0# 0.06fF
C1119 gnd ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C1120 inv_0/in inv_0/op 0.04fF
C1121 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_1/qbar 0.06fF
C1122 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q 0.03fF
C1123 nand_5/a sumffo_1/k 0.02fF
C1124 x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.04fF
C1125 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C1126 vdd inv_1/in 0.30fF
C1127 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/a_10_10# 0.16fF
C1128 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C1129 ffipgarr_0/ffipg_1/ffi_1/qbar vdd 0.33fF
C1130 gnd cla_2/nand_0/w_0_0# 0.01fF
C1131 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C1132 ffipgarr_0/ffi_0/nand_5/w_0_0# vdd 0.10fF
C1133 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C1134 cla_2/nor_1/a_13_6# gnd 0.01fF
C1135 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/b 0.31fF
C1136 clk y1in 0.70fF
C1137 vdd ffo_0/nand_6/w_0_0# 0.10fF
C1138 nand_5/a cla_0/nor_0/a_13_6# 0.01fF
C1139 gnd cla_1/nor_1/w_0_0# 0.01fF
C1140 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_6/w_0_0# 0.06fF
C1141 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.00fF
C1142 inv_9/in nor_4/w_0_0# 0.11fF
C1143 ffo_0/nand_1/a ffo_0/nand_1/w_0_0# 0.06fF
C1144 inv_1/in nand_2/b 0.04fF
C1145 vdd sumffo_3/ffo_0/nand_3/a 0.30fF
C1146 gnd sumffo_1/ffo_0/nand_1/b 0.26fF
C1147 vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C1148 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_0/q 0.73fF
C1149 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C1150 cla_2/inv_0/w_0_6# vdd 0.06fF
C1151 sumffo_1/ffo_0/nand_7/a z2o 0.00fF
C1152 cla_2/p1 gnd 0.69fF
C1153 vdd cla_1/l 0.27fF
C1154 vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.34fF
C1155 gnd sumffo_3/ffo_0/nand_7/a 0.03fF
C1156 sumffo_1/ffo_0/inv_1/w_0_6# sumffo_1/ffo_0/nand_0/b 0.03fF
C1157 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.04fF
C1158 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C1159 ffo_0/inv_0/w_0_6# gnd 0.01fF
C1160 vdd sumffo_3/ffo_0/nand_0/b 0.15fF
C1161 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C1162 inv_5/in cla_0/n 0.13fF
C1163 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_1/q 0.73fF
C1164 ffipgarr_0/ffi_0/nand_2/w_0_0# ffipgarr_0/ffi_0/nand_3/a 0.04fF
C1165 ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd 0.35fF
C1166 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_0/q 0.12fF
C1167 gnd sumffo_1/ffo_0/nand_6/a 0.03fF
C1168 sumffo_2/ffo_0/nand_1/w_0_0# gnd 0.00fF
C1169 cla_2/p0 cla_2/l 0.16fF
C1170 ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd 0.34fF
C1171 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.03fF
C1172 nand_2/b cla_1/l 0.35fF
C1173 inv_5/in nor_3/b 0.04fF
C1174 sumffo_3/k sumffo_3/xor_0/inv_1/op 0.06fF
C1175 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/op 0.04fF
C1176 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C1177 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.31fF
C1178 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C1179 ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 0.13fF
C1180 vdd z1o 0.28fF
C1181 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.06fF
C1182 vdd inv_6/in 0.09fF
C1183 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C1184 inv_7/w_0_6# inv_7/in 0.10fF
C1185 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C1186 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.04fF
C1187 clk ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.13fF
C1188 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C1189 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/d 0.06fF
C1190 gnd ffipgarr_0/ffipg_3/ffi_1/q 0.93fF
C1191 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C1192 vdd sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C1193 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q 0.22fF
C1194 ffipgarr_0/ffipg_0/ffi_0/inv_1/op y1in 0.01fF
C1195 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C1196 gnd sumffo_1/ffo_0/nand_3/b 0.35fF
C1197 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/inv_1/op 0.33fF
C1198 vdd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C1199 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b 0.32fF
C1200 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# vdd 0.10fF
C1201 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q 0.22fF
C1202 clk ffipgarr_0/ffi_0/inv_0/op 0.32fF
C1203 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C1204 cla_1/g0 cla_0/inv_0/op 0.35fF
C1205 clk ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.07fF
C1206 vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.10fF
C1207 gnd cla_0/nor_1/w_0_0# 0.01fF
C1208 vdd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C1209 sumffo_1/k nor_0/a 0.06fF
C1210 gnd sumffo_0/ffo_0/inv_0/op 0.10fF
C1211 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C1212 ffo_0/nand_7/a ffo_0/nand_7/w_0_0# 0.06fF
C1213 vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C1214 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C1215 clk ffo_0/nand_3/b 0.33fF
C1216 vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.10fF
C1217 cla_1/n nor_2/b 0.37fF
C1218 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# vdd 0.10fF
C1219 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C1220 sumffo_2/k cla_1/p0 2.09fF
C1221 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.03fF
C1222 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.04fF
C1223 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.06fF
C1224 cla_0/n sumffo_2/ffo_0/nand_3/b 0.19fF
C1225 clk cla_0/l 0.12fF
C1226 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C1227 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# vdd 0.06fF
C1228 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b 0.13fF
C1229 cla_0/n inv_2/in 0.02fF
C1230 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.06fF
C1231 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# 0.04fF
C1232 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C1233 ffipgarr_0/ffi_0/nand_1/b gnd 0.26fF
C1234 gnd ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.35fF
C1235 sumffo_2/ffo_0/nand_3/a cla_0/l 0.15fF
C1236 vdd x4in 0.04fF
C1237 vdd sumffo_1/ffo_0/nand_7/a 0.30fF
C1238 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.11fF
C1239 inv_7/in vdd 0.34fF
C1240 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C1241 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.04fF
C1242 gnd inv_7/op 0.16fF
C1243 vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.34fF
C1244 clk vdd 12.15fF
C1245 clk ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.06fF
C1246 gnd sumffo_0/ffo_0/nand_3/b 0.35fF
C1247 ffo_0/nand_0/b ffo_0/nand_2/w_0_0# 0.06fF
C1248 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C1249 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# 0.04fF
C1250 z3o sumffo_2/ffo_0/nand_6/a 0.31fF
C1251 gnd ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.26fF
C1252 inv_4/op sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C1253 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C1254 vdd sumffo_2/ffo_0/nand_3/a 0.30fF
C1255 cla_0/n inv_3/w_0_6# 0.00fF
C1256 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C1257 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C1258 couto ffo_0/qbar 0.32fF
C1259 ffipgarr_0/ffi_0/inv_1/op cinin 0.01fF
C1260 cla_1/p0 cla_2/p0 0.24fF
C1261 vdd sumffo_2/ffo_0/nand_1/b 0.31fF
C1262 vdd inv_0/op 0.17fF
C1263 sumffo_1/xor_0/w_n3_4# sumffo_1/ffo_0/d 0.02fF
C1264 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C1265 gnd ffipgarr_0/ffipg_3/ffi_1/qbar 0.34fF
C1266 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in 0.04fF
C1267 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C1268 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.31fF
C1269 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.06fF
C1270 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C1271 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C1272 vdd ffo_0/qbar 0.28fF
C1273 inv_3/in nor_2/b 0.04fF
C1274 ffipgarr_0/ffi_0/nand_7/a gnd 0.03fF
C1275 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/q 0.31fF
C1276 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.04fF
C1277 gnd cla_1/inv_0/in 0.35fF
C1278 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_1/w_0_6# 0.03fF
C1279 sumffo_0/ffo_0/nand_7/a sumffo_0/sbar 0.31fF
C1280 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C1281 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.06fF
C1282 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.20fF
C1283 ffo_0/nand_3/a vdd 0.30fF
C1284 vdd sumffo_1/ffo_0/d 0.04fF
C1285 sumffo_2/ffo_0/nand_0/b gnd 0.38fF
C1286 cla_2/inv_0/op cla_2/nand_0/w_0_0# 0.06fF
C1287 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.03fF
C1288 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.13fF
C1289 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.06fF
C1290 vdd ffipgarr_0/ffipg_1/ffi_0/qbar 0.33fF
C1291 cla_1/inv_0/op cla_2/g0 0.35fF
C1292 clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C1293 ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd 0.17fF
C1294 ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd 1.63fF
C1295 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C1296 vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.34fF
C1297 gnd cla_2/inv_0/op 0.10fF
C1298 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.06fF
C1299 ffo_0/d ffo_0/nand_2/w_0_0# 0.06fF
C1300 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C1301 vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C1302 vdd ffipgarr_0/ffipg_2/ffi_0/q 0.38fF
C1303 cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C1304 ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd 1.63fF
C1305 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.31fF
C1306 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a 0.00fF
C1307 clk ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C1308 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C1309 gnd cla_1/nand_0/w_0_0# 0.01fF
C1310 vdd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C1311 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C1312 gnd sumffo_0/k 0.41fF
C1313 nand_5/a ffipgarr_0/ffi_0/nand_6/a 0.31fF
C1314 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.30fF
C1315 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# vdd 0.06fF
C1316 nor_0/b inv_0/in 0.16fF
C1317 z1o sumffo_0/ffo_0/nand_6/a 0.31fF
C1318 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q 0.32fF
C1319 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.04fF
C1320 sumffo_2/ffo_0/nand_1/a_13_n26# gnd 0.01fF
C1321 sumffo_3/ffo_0/nand_6/a sumffo_3/sbar 0.00fF
C1322 clk sumffo_0/ffo_0/nand_1/b 0.45fF
C1323 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_1/op 0.52fF
C1324 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.31fF
C1325 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.00fF
C1326 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C1327 gnd ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.03fF
C1328 vdd z3o 0.28fF
C1329 vdd sumffo_2/ffo_0/nand_4/w_0_0# 0.10fF
C1330 clk ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.07fF
C1331 vdd sumffo_1/ffo_0/nand_0/b 0.15fF
C1332 vdd sumffo_0/ffo_0/nand_1/w_0_0# 0.10fF
C1333 sumffo_1/sbar gnd 0.34fF
C1334 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C1335 gnd ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.03fF
C1336 sumffo_0/ffo_0/nand_7/w_0_0# vdd 0.10fF
C1337 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.31fF
C1338 vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.17fF
C1339 nor_3/w_0_0# nor_3/b 0.06fF
C1340 gnd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.00fF
C1341 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.04fF
C1342 nor_4/b nor_4/w_0_0# 0.06fF
C1343 sumffo_3/ffo_0/nand_2/w_0_0# vdd 0.10fF
C1344 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C1345 vdd sumffo_1/ffo_0/nand_1/w_0_0# 0.10fF
C1346 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1347 inv_7/w_0_6# cla_2/l 0.06fF
C1348 nand_5/a gnd 0.91fF
C1349 sumffo_2/ffo_0/nand_1/a cla_0/l 0.15fF
C1350 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_0/op 0.08fF
C1351 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.07fF
C1352 vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.17fF
C1353 inv_0/op nand_0/w_0_0# 0.06fF
C1354 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C1355 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q 0.29fF
C1356 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a 0.00fF
C1357 cla_2/nor_0/w_0_0# cla_2/p0 0.06fF
C1358 ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd 0.39fF
C1359 vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.10fF
C1360 gnd ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.35fF
C1361 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C1362 gnd ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# 0.01fF
C1363 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b 0.13fF
C1364 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1365 gnd sumffo_2/xor_0/inv_0/op 0.17fF
C1366 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.06fF
C1367 inv_3/w_0_6# cla_1/l 0.06fF
C1368 clk ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.06fF
C1369 vdd sumffo_2/ffo_0/nand_1/a 0.30fF
C1370 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.06fF
C1371 clk sumffo_0/ffo_0/nand_6/a 0.13fF
C1372 clk x3in 0.70fF
C1373 cla_0/n gnd 0.52fF
C1374 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C1375 vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.10fF
C1376 vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.17fF
C1377 clk ffipgarr_0/ffi_0/nand_3/a 0.13fF
C1378 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.13fF
C1379 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C1380 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.31fF
C1381 nor_0/b ffipgarr_0/ffipg_0/ffi_1/q 1.27fF
C1382 nor_0/b ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C1383 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q 0.32fF
C1384 cla_2/l cla_0/l 0.40fF
C1385 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.75fF
C1386 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_6/w_0_0# 0.06fF
C1387 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C1388 sumffo_1/ffo_0/inv_0/w_0_6# sumffo_1/ffo_0/d 0.06fF
C1389 sumffo_2/sbar vdd 0.28fF
C1390 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.00fF
C1391 nor_3/b gnd 0.10fF
C1392 inv_8/w_0_6# vdd 0.15fF
C1393 ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd 0.03fF
C1394 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C1395 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b 0.13fF
C1396 vdd sumffo_0/ffo_0/nand_0/b 0.15fF
C1397 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C1398 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# vdd 0.11fF
C1399 vdd cla_2/l 0.40fF
C1400 cla_0/n sumffo_2/ffo_0/nand_1/w_0_0# 0.13fF
C1401 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C1402 vdd cla_1/inv_0/op 0.17fF
C1403 gnd ffo_0/nand_1/b 0.26fF
C1404 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/w_0_0# 0.06fF
C1405 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.31fF
C1406 vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.10fF
C1407 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1408 inv_4/op sumffo_3/xor_0/inv_1/op 0.22fF
C1409 vdd sumffo_3/ffo_0/nand_4/w_0_0# 0.10fF
C1410 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/ffi_0/nand_0/w_0_0# 0.06fF
C1411 clk y3in 0.70fF
C1412 gnd ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.03fF
C1413 vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.34fF
C1414 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C1415 vdd sumffo_0/ffo_0/nand_0/w_0_0# 0.10fF
C1416 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1417 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C1418 gnd cla_1/g0 0.76fF
C1419 clk sumffo_2/ffo_0/nand_3/b 0.33fF
C1420 ffipgarr_0/ffipg_2/ffi_1/inv_1/op x3in 0.01fF
C1421 vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C1422 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C1423 ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd 0.34fF
C1424 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1425 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C1426 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C1427 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C1428 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.30fF
C1429 gnd nor_0/a 0.29fF
C1430 ffo_0/nand_0/b ffo_0/nand_1/a 0.13fF
C1431 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_3/b 0.31fF
C1432 ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd 0.39fF
C1433 gnd ffipgarr_0/ffipg_0/ffi_1/qbar 0.34fF
C1434 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C1435 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.06fF
C1436 cla_0/n nor_1/w_0_0# 0.06fF
C1437 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b 0.32fF
C1438 sumffo_0/ffo_0/nand_1/a gnd 0.03fF
C1439 vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C1440 nand_5/a inv_7/op 0.38fF
C1441 sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/inv_0/op 0.08fF
C1442 vdd sumffo_1/ffo_0/inv_0/op 0.17fF
C1443 gnd sumffo_0/xor_0/inv_0/op 0.17fF
C1444 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# x3in 0.06fF
C1445 vdd ffo_0/nand_2/w_0_0# 0.10fF
C1446 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C1447 gnd sumffo_3/ffo_0/inv_0/op 0.32fF
C1448 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C1449 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.30fF
C1450 nor_0/b vdd 0.90fF
C1451 vdd ffipgarr_0/ffi_0/nand_0/w_0_0# 0.10fF
C1452 clk ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.32fF
C1453 inv_1/in gnd 0.22fF
C1454 vdd sumffo_2/ffo_0/nand_6/w_0_0# 0.10fF
C1455 vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# 0.10fF
C1456 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.32fF
C1457 ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 1.40fF
C1458 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C1459 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_0/q 0.12fF
C1460 ffipgarr_0/ffipg_1/ffi_1/qbar gnd 0.34fF
C1461 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.06fF
C1462 cla_1/p0 cla_0/l 0.02fF
C1463 couto ffo_0/nand_6/a 0.31fF
C1464 nor_3/w_0_0# inv_6/in 0.11fF
C1465 vdd sumffo_3/xor_0/inv_1/op 0.15fF
C1466 cla_2/g0 cla_2/nor_1/w_0_0# 0.06fF
C1467 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.33fF
C1468 ffipgarr_0/ffi_0/nand_6/w_0_0# vdd 0.10fF
C1469 nor_1/b cla_0/l 0.10fF
C1470 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.04fF
C1471 vdd cla_0/g0 0.50fF
C1472 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# vdd 0.11fF
C1473 clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.13fF
C1474 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C1475 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C1476 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/q 0.31fF
C1477 ffipgarr_0/ffi_0/nand_7/a nand_5/a 0.00fF
C1478 ffipgarr_0/ffi_0/nand_1/a clk 0.13fF
C1479 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C1480 z4o sumffo_3/sbar 0.32fF
C1481 gnd sumffo_3/ffo_0/nand_3/a 0.03fF
C1482 vdd cla_1/p0 0.44fF
C1483 vdd ffo_0/nand_6/a 0.30fF
C1484 x3in ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.04fF
C1485 gnd cla_1/l 0.18fF
C1486 x1in ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C1487 cla_1/n nor_2/w_0_0# 0.06fF
C1488 gnd ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.03fF
C1489 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.04fF
C1490 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.04fF
C1491 x2in ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.01fF
C1492 vdd nor_1/b 0.35fF
C1493 gnd sumffo_3/ffo_0/nand_0/b 0.38fF
C1494 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C1495 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1496 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1497 nand_2/b cla_0/g0 1.01fF
C1498 sumffo_1/ffo_0/nand_2/w_0_0# sumffo_1/ffo_0/d 0.06fF
C1499 sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# 0.02fF
C1500 cla_1/n cla_2/g0 0.13fF
C1501 clk ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1502 cla_1/p0 nand_2/b 2.00fF
C1503 ffipgarr_0/ffipg_3/ffi_0/nand_3/a clk 0.13fF
C1504 ffo_0/nand_0/b ffo_0/inv_0/op 0.32fF
C1505 ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd 1.63fF
C1506 sumffo_2/ffo_0/nand_4/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C1507 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.30fF
C1508 vdd sumffo_3/ffo_0/nand_6/a 0.30fF
C1509 ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd 0.03fF
C1510 vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.34fF
C1511 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/q 0.00fF
C1512 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C1513 nand_5/a sumffo_0/k 0.41fF
C1514 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C1515 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.06fF
C1516 gnd ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.26fF
C1517 ffipgarr_0/ffi_0/inv_1/w_0_6# clk 0.06fF
C1518 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C1519 z1o gnd 0.52fF
C1520 gnd inv_6/in 0.24fF
C1521 clk ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.06fF
C1522 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b 0.31fF
C1523 inv_5/in cla_2/l 0.03fF
C1524 clk ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1525 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C1526 x2in vdd 0.04fF
C1527 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.04fF
C1528 cla_0/n cla_1/nand_0/w_0_0# 0.01fF
C1529 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.31fF
C1530 vdd y2in 0.04fF
C1531 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C1532 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C1533 vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.10fF
C1534 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C1535 y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1536 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1537 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1538 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.03fF
C1539 ffipgarr_0/ffipg_2/ffi_0/inv_0/op ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.06fF
C1540 vdd cla_0/inv_0/w_0_6# 0.06fF
C1541 sumffo_3/ffo_0/nand_0/w_0_0# vdd 0.10fF
C1542 ffipgarr_0/ffipg_2/ffi_0/nand_1/b vdd 0.31fF
C1543 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.13fF
C1544 cla_1/g0 cla_1/inv_0/in 0.16fF
C1545 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q 0.32fF
C1546 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.04fF
C1547 cla_0/nand_0/w_0_0# cla_0/l 0.15fF
C1548 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_3/b 0.00fF
C1549 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C1550 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1551 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.06fF
C1552 ffo_0/d ffo_0/inv_0/op 0.04fF
C1553 vdd sumffo_0/ffo_0/nand_7/a 0.30fF
C1554 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.31fF
C1555 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/q 0.31fF
C1556 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C1557 sumffo_1/ffo_0/nand_6/w_0_0# sumffo_1/ffo_0/nand_6/a 0.06fF
C1558 sumffo_0/ffo_0/d sumffo_0/xor_0/a_10_10# 0.45fF
C1559 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.03fF
C1560 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C1561 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C1562 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.00fF
C1563 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar 0.32fF
C1564 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C1565 gnd x4in 0.19fF
C1566 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.13fF
C1567 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.32fF
C1568 gnd sumffo_1/ffo_0/nand_7/a 0.03fF
C1569 cla_0/g0 nand_0/w_0_0# 0.06fF
C1570 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b 0.13fF
C1571 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C1572 ffipgarr_0/ffi_0/nand_3/b vdd 0.39fF
C1573 vdd cla_0/nand_0/w_0_0# 0.10fF
C1574 inv_7/in gnd 0.13fF
C1575 vdd sumffo_2/ffo_0/nand_3/w_0_0# 0.11fF
C1576 gnd ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.03fF
C1577 clk gnd 8.12fF
C1578 clk sumffo_1/ffo_0/nand_1/b 0.45fF
C1579 gnd cla_1/nor_1/a_13_6# 0.01fF
C1580 ffo_0/nand_7/a couto 0.00fF
C1581 vdd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C1582 sumffo_1/k cla_0/g0 0.07fF
C1583 vdd cla_2/nor_0/w_0_0# 0.31fF
C1584 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1585 gnd sumffo_2/ffo_0/nand_3/a 0.03fF
C1586 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C1587 vdd cla_2/nor_1/w_0_0# 0.31fF
C1588 cinin ffipgarr_0/ffi_0/inv_0/op 0.04fF
C1589 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.11fF
C1590 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.04fF
C1591 sumffo_1/k cla_1/p0 0.05fF
C1592 cla_0/nand_0/w_0_0# nand_2/b 0.01fF
C1593 vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.10fF
C1594 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C1595 nor_2/w_0_0# nor_2/b 0.06fF
C1596 gnd inv_0/op 0.10fF
C1597 gnd sumffo_2/ffo_0/nand_1/b 0.38fF
C1598 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C1599 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# 0.04fF
C1600 vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C1601 sumffo_0/k nor_0/a 0.05fF
C1602 cla_1/n cla_0/l 0.18fF
C1603 ffo_0/nand_7/a vdd 0.30fF
C1604 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1605 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C1606 clk sumffo_1/ffo_0/nand_6/a 0.13fF
C1607 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C1608 vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.10fF
C1609 gnd ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.26fF
C1610 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C1611 sumffo_3/k cla_2/p0 0.09fF
C1612 inv_2/op sumffo_2/k 0.09fF
C1613 gnd ffo_0/qbar 0.34fF
C1614 ffo_0/nand_1/a ffo_0/nand_3/b 0.00fF
C1615 sumffo_0/xor_0/inv_0/op sumffo_0/k 0.27fF
C1616 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.06fF
C1617 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1618 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.04fF
C1619 nor_4/b inv_8/w_0_6# 0.03fF
C1620 ffo_0/nand_3/a gnd 0.14fF
C1621 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C1622 gnd sumffo_1/ffo_0/d 0.37fF
C1623 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_0/ffi_1/qbar 0.04fF
C1624 cla_1/n vdd 0.28fF
C1625 sumffo_3/k sumffo_3/xor_0/inv_0/op 0.27fF
C1626 sumffo_2/xor_0/w_n3_4# sumffo_2/xor_0/inv_1/op 0.06fF
C1627 vdd cla_0/inv_0/in 0.05fF
C1628 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.31fF
C1629 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.00fF
C1630 gnd ffipgarr_0/ffipg_1/ffi_0/qbar 0.34fF
C1631 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C1632 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.31fF
C1633 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C1634 vdd sumffo_1/ffo_0/nand_3/a 0.30fF
C1635 ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd 0.10fF
C1636 clk sumffo_1/ffo_0/nand_3/b 0.33fF
C1637 ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd 0.22fF
C1638 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.75fF
C1639 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C1640 gnd ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.03fF
C1641 vdd ffo_0/nand_1/w_0_0# 0.10fF
C1642 sumffo_2/k cla_2/p0 0.05fF
C1643 sumffo_2/ffo_0/nand_7/w_0_0# z3o 0.04fF
C1644 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C1645 vdd cinin 0.04fF
C1646 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# y3in 0.06fF
C1647 gnd ffipgarr_0/ffipg_2/ffi_0/q 2.62fF
C1648 ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd 0.22fF
C1649 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.11fF
C1650 nand_5/a nor_0/a 0.26fF
C1651 ffo_0/nand_1/a vdd 0.30fF
C1652 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a 0.13fF
C1653 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.00fF
C1654 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C1655 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.30fF
C1656 sumffo_1/xor_0/inv_1/op vdd 0.15fF
C1657 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C1658 inv_0/in nor_0/w_0_0# 0.11fF
C1659 vdd sumffo_2/ffo_0/d 0.04fF
C1660 gnd ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.14fF
C1661 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/d 0.06fF
C1662 cla_0/n cla_1/g0 0.13fF
C1663 vdd sumffo_2/ffo_0/nand_7/a 0.30fF
C1664 nand_5/a sumffo_0/xor_0/inv_0/op 0.20fF
C1665 clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.13fF
C1666 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.31fF
C1667 vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1668 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# gnd 0.01fF
C1669 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# sumffo_3/k 0.45fF
C1670 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1671 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C1672 inv_3/in cla_0/l 0.06fF
C1673 cla_0/n sumffo_2/ffo_0/nand_2/w_0_0# 0.13fF
C1674 gnd z3o 0.52fF
C1675 vdd sumffo_2/ffo_0/inv_0/op 0.17fF
C1676 gnd sumffo_1/ffo_0/nand_0/b 0.45fF
C1677 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.30fF
C1678 cla_0/inv_0/w_0_6# cla_0/inv_0/op 0.03fF
C1679 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C1680 nand_5/a inv_1/in 0.13fF
C1681 sumffo_1/xor_0/inv_1/op nand_2/b 0.22fF
C1682 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op 1.63fF
C1683 inv_7/in inv_7/op 0.04fF
C1684 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.04fF
C1685 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/q 0.31fF
C1686 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C1687 vdd z4o 0.28fF
C1688 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.31fF
C1689 gnd ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.10fF
C1690 cla_0/l inv_1/w_0_6# 0.28fF
C1691 clk sumffo_0/ffo_0/nand_3/b 0.33fF
C1692 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.31fF
C1693 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.04fF
C1694 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C1695 ffipgarr_0/ffipg_2/ffi_0/inv_1/op y3in 0.01fF
C1696 inv_3/in vdd 0.30fF
C1697 ffo_0/nand_1/b ffo_0/nand_5/w_0_0# 0.06fF
C1698 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_1/ffi_1/q 0.06fF
C1699 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.06fF
C1700 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C1701 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C1702 vdd sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1703 nor_1/b inv_2/in 0.16fF
C1704 vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C1705 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C1706 gnd ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.10fF
C1707 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1708 vdd inv_1/w_0_6# 0.15fF
C1709 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C1710 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# 0.04fF
C1711 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.10fF
C1712 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# vdd 0.06fF
C1713 sumffo_2/sbar sumffo_2/ffo_0/nand_7/w_0_0# 0.06fF
C1714 ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd 0.35fF
C1715 clk ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.06fF
C1716 vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.10fF
C1717 inv_3/in nand_2/b 0.13fF
C1718 cla_1/p0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C1719 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.06fF
C1720 clk sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C1721 inv_2/op sumffo_2/xor_0/a_10_10# 0.12fF
C1722 gnd sumffo_2/ffo_0/nand_1/a 0.06fF
C1723 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C1724 ffipgarr_0/ffipg_2/ffi_1/q sumffo_2/k 2.17fF
C1725 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# y2in 0.06fF
C1726 vdd ffo_0/inv_0/op 0.17fF
C1727 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.04fF
C1728 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a 0.31fF
C1729 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.06fF
C1730 nand_2/b inv_1/w_0_6# 0.01fF
C1731 clk sumffo_2/ffo_0/nand_0/b 0.04fF
C1732 gnd ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.34fF
C1733 sumffo_3/k cla_2/g0 0.10fF
C1734 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.33fF
C1735 vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.17fF
C1736 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C1737 z1o sumffo_0/ffo_0/nand_6/w_0_0# 0.06fF
C1738 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.06fF
C1739 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C1740 vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.34fF
C1741 couto ffo_0/nand_7/w_0_0# 0.04fF
C1742 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C1743 sumffo_2/sbar gnd 0.34fF
C1744 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C1745 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C1746 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.33fF
C1747 sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# 0.04fF
C1748 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C1749 vdd nor_2/b 0.35fF
C1750 ffipgarr_0/ffipg_2/ffi_1/nand_1/b vdd 0.31fF
C1751 vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.10fF
C1752 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar 0.32fF
C1753 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.27fF
C1754 cla_0/g0 ffipgarr_0/ffipg_1/ffi_1/q 0.84fF
C1755 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C1756 gnd sumffo_0/ffo_0/nand_0/b 0.38fF
C1757 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.04fF
C1758 inv_4/in cla_1/n 0.02fF
C1759 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_3/b 0.04fF
C1760 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.45fF
C1761 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.30fF
C1762 ffo_0/nand_7/w_0_0# vdd 0.12fF
C1763 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1764 sumffo_2/ffo_0/nand_1/w_0_0# sumffo_2/ffo_0/nand_1/a 0.06fF
C1765 cla_1/p0 ffipgarr_0/ffipg_1/ffi_1/q 0.22fF
C1766 gnd cla_2/l 0.36fF
C1767 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C1768 cla_2/p1 cla_2/l 0.02fF
C1769 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C1770 gnd cla_1/inv_0/op 0.15fF
C1771 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C1772 vdd ffipgarr_0/ffipg_0/ffi_0/qbar 0.33fF
C1773 gnd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.00fF
C1774 vdd sumffo_0/xor_0/w_n3_4# 0.12fF
C1775 ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 0.22fF
C1776 vdd ffipgarr_0/ffi_0/inv_1/op 1.67fF
C1777 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C1778 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C1779 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q 0.21fF
C1780 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C1781 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C1782 nor_0/b ffipgarr_0/ffi_0/nand_6/a 0.00fF
C1783 gnd ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.03fF
C1784 clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.13fF
C1785 sumffo_1/xor_0/inv_1/op sumffo_1/k 0.06fF
C1786 sumffo_1/sbar sumffo_1/ffo_0/nand_7/a 0.31fF
C1787 gnd cla_0/nor_1/a_13_6# 0.01fF
C1788 sumffo_3/k sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C1789 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_6/w_0_0# 0.06fF
C1790 vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.17fF
C1791 sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d 0.06fF
C1792 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/b 0.06fF
C1793 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C1794 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.30fF
C1795 nor_3/b inv_6/in 0.16fF
C1796 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# 0.04fF
C1797 ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd 0.03fF
C1798 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.13fF
C1799 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# cla_0/g0 0.04fF
C1800 vdd inv_8/in 0.30fF
C1801 gnd ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.14fF
C1802 inv_9/in Gnd 0.23fF
C1803 nor_4/w_0_0# Gnd 1.81fF
C1804 nor_4/b Gnd 0.81fF
C1805 inv_8/in Gnd 0.22fF
C1806 inv_8/w_0_6# Gnd 1.40fF
C1807 inv_7/in Gnd 0.22fF
C1808 inv_7/w_0_6# Gnd 1.40fF
C1809 nor_4/a Gnd 0.27fF
C1810 nor_3/b Gnd 0.54fF
C1811 inv_5/in Gnd 0.22fF
C1812 inv_5/w_0_6# Gnd 1.40fF
C1813 cla_2/n Gnd 0.32fF
C1814 inv_6/in Gnd 0.23fF
C1815 nor_3/w_0_0# Gnd 1.81fF
C1816 nor_2/b Gnd 0.92fF
C1817 cla_1/n Gnd 0.20fF
C1818 inv_4/in Gnd 0.23fF
C1819 nor_2/w_0_0# Gnd 1.81fF
C1820 cla_0/n Gnd 0.68fF
C1821 inv_3/in Gnd 0.22fF
C1822 inv_3/w_0_6# Gnd 1.40fF
C1823 inv_2/op Gnd 1.94fF
C1824 inv_2/in Gnd 0.23fF
C1825 nor_1/w_0_0# Gnd 1.81fF
C1826 nor_1/b Gnd 0.85fF
C1827 inv_1/in Gnd 0.22fF
C1828 inv_1/w_0_6# Gnd 1.40fF
C1829 inv_0/in Gnd 0.23fF
C1830 nor_0/w_0_0# Gnd 1.81fF
C1831 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1832 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1833 ffo_0/nand_7/a Gnd 0.30fF
C1834 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1835 ffo_0/qbar Gnd 0.42fF
C1836 ffo_0/nand_6/a Gnd 0.30fF
C1837 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1838 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1839 ffo_0/nand_3/b Gnd 0.43fF
C1840 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1841 ffo_0/nand_3/a Gnd 0.30fF
C1842 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1843 ffo_0/nand_0/b Gnd 0.63fF
C1844 ffo_0/d Gnd 0.60fF
C1845 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1846 ffo_0/inv_0/op Gnd 0.26fF
C1847 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1848 ffo_0/nand_1/a Gnd 0.30fF
C1849 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1850 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1851 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1852 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1853 inv_4/op Gnd 1.54fF
C1854 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1855 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1856 sumffo_3/k Gnd 3.28fF
C1857 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1858 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1859 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1860 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1861 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1862 sumffo_3/sbar Gnd 0.43fF
C1863 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1864 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1865 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1866 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1867 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1868 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1869 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1870 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1871 sumffo_3/ffo_0/d Gnd 0.64fF
C1872 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1873 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1874 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1875 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1876 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1877 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1878 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1879 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1880 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1881 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1882 sumffo_1/k Gnd 2.61fF
C1883 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1884 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1885 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1886 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1887 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1888 sumffo_1/sbar Gnd 0.43fF
C1889 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1890 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1891 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1892 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1893 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1894 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1895 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1896 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1897 sumffo_1/ffo_0/d Gnd 0.64fF
C1898 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1899 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1900 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1901 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1902 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1903 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1904 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1905 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1906 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1907 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1908 sumffo_2/k Gnd 1.72fF
C1909 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1910 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1911 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1912 gnd Gnd 47.57fF
C1913 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1914 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1915 sumffo_2/sbar Gnd 0.43fF
C1916 vdd Gnd 26.61fF
C1917 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1918 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1919 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1920 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1921 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1922 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1923 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1924 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1925 sumffo_2/ffo_0/d Gnd 0.64fF
C1926 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1927 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1928 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1929 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1930 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1931 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1932 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1933 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1934 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1935 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1936 sumffo_0/k Gnd 3.08fF
C1937 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1938 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1939 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1940 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1941 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1942 sumffo_0/sbar Gnd 0.43fF
C1943 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1944 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1945 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1946 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1947 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1948 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1949 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1950 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1951 sumffo_0/ffo_0/d Gnd 0.64fF
C1952 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1953 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1954 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1955 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1956 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1957 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1958 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1959 cla_2/inv_0/in Gnd 0.27fF
C1960 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1961 cla_2/inv_0/op Gnd 0.26fF
C1962 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1963 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1964 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1965 ffipgarr_0/ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1966 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1967 ffipgarr_0/ffipg_3/ffi_1/qbar Gnd 0.42fF
C1968 ffipgarr_0/ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1969 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1970 ffipgarr_0/ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1971 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1972 ffipgarr_0/ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1973 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1974 ffipgarr_0/ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1975 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1976 x4in Gnd 0.52fF
C1977 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1978 ffipgarr_0/ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1979 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1980 ffipgarr_0/ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1981 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1982 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1983 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1984 ffipgarr_0/ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1985 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1986 ffipgarr_0/ffipg_3/ffi_0/qbar Gnd 0.42fF
C1987 ffipgarr_0/ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1988 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1989 ffipgarr_0/ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1990 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1991 ffipgarr_0/ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1992 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1993 ffipgarr_0/ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1994 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1995 y4in Gnd 0.52fF
C1996 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1997 ffipgarr_0/ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1998 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C1999 ffipgarr_0/ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C2000 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2001 cla_2/p1 Gnd 0.89fF
C2002 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2003 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2004 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2005 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2006 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2007 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2008 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2009 cla_2/g1 Gnd 0.66fF
C2010 ffipgarr_0/ffipg_3/ffi_0/q Gnd 2.68fF
C2011 ffipgarr_0/ffipg_3/ffi_1/q Gnd 2.93fF
C2012 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2013 ffipgarr_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2014 ffipgarr_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2015 ffipgarr_0/ffi_0/nand_7/a Gnd 0.30fF
C2016 ffipgarr_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2017 nor_0/b Gnd 1.09fF
C2018 ffipgarr_0/ffi_0/nand_6/a Gnd 0.30fF
C2019 ffipgarr_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2020 ffipgarr_0/ffi_0/inv_1/op Gnd 0.89fF
C2021 ffipgarr_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2022 ffipgarr_0/ffi_0/nand_3/b Gnd 0.43fF
C2023 ffipgarr_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2024 ffipgarr_0/ffi_0/nand_3/a Gnd 0.30fF
C2025 ffipgarr_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2026 clk Gnd 17.25fF
C2027 cinin Gnd 0.52fF
C2028 ffipgarr_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2029 ffipgarr_0/ffi_0/inv_0/op Gnd 0.26fF
C2030 ffipgarr_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2031 ffipgarr_0/ffi_0/nand_1/a Gnd 0.30fF
C2032 ffipgarr_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2033 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2034 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2035 ffipgarr_0/ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C2036 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2037 ffipgarr_0/ffipg_2/ffi_1/qbar Gnd 0.42fF
C2038 ffipgarr_0/ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C2039 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2040 ffipgarr_0/ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C2041 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2042 ffipgarr_0/ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C2043 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2044 ffipgarr_0/ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C2045 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2046 x3in Gnd 0.52fF
C2047 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2048 ffipgarr_0/ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C2049 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2050 ffipgarr_0/ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C2051 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2052 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2053 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2054 ffipgarr_0/ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C2055 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2056 ffipgarr_0/ffipg_2/ffi_0/qbar Gnd 0.42fF
C2057 ffipgarr_0/ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C2058 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2059 ffipgarr_0/ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C2060 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2061 ffipgarr_0/ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C2062 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2063 ffipgarr_0/ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C2064 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2065 y3in Gnd 0.52fF
C2066 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2067 ffipgarr_0/ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C2068 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2069 ffipgarr_0/ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C2070 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2071 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2072 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2073 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2074 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2075 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2076 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2077 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2078 ffipgarr_0/ffipg_2/ffi_0/q Gnd 2.68fF
C2079 ffipgarr_0/ffipg_2/ffi_1/q Gnd 2.93fF
C2080 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2081 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2082 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2083 ffipgarr_0/ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C2084 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2085 ffipgarr_0/ffipg_1/ffi_1/qbar Gnd 0.42fF
C2086 ffipgarr_0/ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C2087 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2088 ffipgarr_0/ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C2089 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2090 ffipgarr_0/ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C2091 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2092 ffipgarr_0/ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C2093 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2094 x2in Gnd 0.52fF
C2095 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2096 ffipgarr_0/ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C2097 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2098 ffipgarr_0/ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C2099 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2100 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2101 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2102 ffipgarr_0/ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C2103 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2104 ffipgarr_0/ffipg_1/ffi_0/qbar Gnd 0.42fF
C2105 ffipgarr_0/ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C2106 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2107 ffipgarr_0/ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C2108 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2109 ffipgarr_0/ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C2110 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2111 ffipgarr_0/ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C2112 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2113 y2in Gnd 0.43fF
C2114 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2115 ffipgarr_0/ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C2116 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2117 ffipgarr_0/ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C2118 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2119 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2120 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2121 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2122 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2123 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2124 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2125 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2126 ffipgarr_0/ffipg_1/ffi_0/q Gnd 2.68fF
C2127 ffipgarr_0/ffipg_1/ffi_1/q Gnd 2.93fF
C2128 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2129 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2130 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2131 ffipgarr_0/ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C2132 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2133 ffipgarr_0/ffipg_0/ffi_1/qbar Gnd 0.42fF
C2134 ffipgarr_0/ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C2135 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2136 ffipgarr_0/ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C2137 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2138 ffipgarr_0/ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C2139 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2140 ffipgarr_0/ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C2141 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2142 x1in Gnd 0.42fF
C2143 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2144 ffipgarr_0/ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C2145 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2146 ffipgarr_0/ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C2147 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2148 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2149 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2150 ffipgarr_0/ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C2151 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2152 ffipgarr_0/ffipg_0/ffi_0/qbar Gnd 0.42fF
C2153 ffipgarr_0/ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C2154 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2155 ffipgarr_0/ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C2156 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2157 ffipgarr_0/ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C2158 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2159 ffipgarr_0/ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C2160 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2161 y1in Gnd 0.52fF
C2162 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2163 ffipgarr_0/ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C2164 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2165 ffipgarr_0/ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C2166 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2167 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2168 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2169 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2170 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2171 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2172 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2173 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2174 ffipgarr_0/ffipg_0/ffi_0/q Gnd 2.68fF
C2175 ffipgarr_0/ffipg_0/ffi_1/q Gnd 2.93fF
C2176 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2177 cla_2/p0 Gnd 1.30fF
C2178 cla_1/nor_1/w_0_0# Gnd 1.23fF
C2179 cla_1/l Gnd 0.31fF
C2180 cla_1/nor_0/w_0_0# Gnd 1.23fF
C2181 cla_1/inv_0/in Gnd 0.27fF
C2182 cla_1/inv_0/w_0_6# Gnd 0.58fF
C2183 cla_1/inv_0/op Gnd 0.26fF
C2184 cla_1/nand_0/w_0_0# Gnd 0.82fF
C2185 inv_7/op Gnd 0.30fF
C2186 cla_0/nor_1/w_0_0# Gnd 1.23fF
C2187 cla_0/l Gnd 7.26fF
C2188 cla_0/nor_0/w_0_0# Gnd 1.23fF
C2189 cla_0/inv_0/in Gnd 0.27fF
C2190 cla_0/inv_0/w_0_6# Gnd 0.58fF
C2191 cla_1/g0 Gnd 2.32fF
C2192 cla_0/inv_0/op Gnd 0.26fF
C2193 cla_0/nand_0/w_0_0# Gnd 0.82fF
C2194 cla_2/l Gnd 1.11fF
C2195 nand_2/b Gnd 0.27fF
C2196 inv_0/op Gnd 0.26fF
C2197 nand_0/w_0_0# Gnd 0.82fF
