magic
tech scmos
timestamp 1619188927
<< metal1 >>
rect -3 1270 97 1273
rect 102 1270 546 1273
rect 3 1263 410 1266
rect 3 1256 6 1263
rect -3 1252 0 1255
rect 241 1212 260 1215
rect 241 1156 254 1159
rect -3 1153 0 1156
rect -3 1083 0 1086
rect 251 1047 254 1156
rect 257 1056 260 1212
rect 278 1145 293 1148
rect 278 1054 281 1145
rect 415 1143 418 1146
rect 641 1137 644 1140
rect 262 1051 281 1054
rect 251 1044 497 1047
rect 479 1014 484 1019
rect 494 998 497 1044
rect 539 1026 542 1036
rect 563 1023 572 1026
rect 970 1001 971 1004
rect 494 995 505 998
rect 563 994 572 997
rect 606 993 612 996
rect 617 993 618 996
rect 490 989 505 992
rect 566 988 572 991
rect 539 975 542 978
rect 566 966 569 988
rect 495 963 569 966
rect 572 963 576 966
rect 611 939 618 942
rect -3 876 0 879
rect 611 874 614 939
rect 481 871 614 874
rect -3 802 0 805
rect 481 738 484 871
rect 606 762 609 775
rect 568 748 572 751
rect 479 735 484 738
rect 567 742 572 745
rect 630 743 633 746
rect 505 732 509 735
rect 567 734 570 742
rect 563 729 570 734
rect 636 727 643 730
rect 12 718 17 721
rect 636 717 639 727
rect 677 717 680 730
rect 630 714 639 717
rect 606 713 630 714
rect 490 708 507 711
rect 1077 693 1080 696
rect 638 686 643 689
rect 701 685 725 688
rect 853 687 854 690
rect 487 674 490 682
rect 501 680 507 683
rect 628 682 643 683
rect 633 680 643 682
rect 487 671 507 674
rect 640 654 643 664
rect 677 661 680 669
rect 627 651 643 654
rect -3 595 0 598
rect 722 551 725 634
rect 480 548 725 551
rect -3 521 0 524
rect 480 457 483 548
rect 617 481 620 494
rect 579 467 583 470
rect 578 461 583 464
rect 641 462 644 465
rect 508 451 520 454
rect 578 453 581 461
rect 574 448 581 453
rect 647 446 654 449
rect 647 436 650 446
rect 688 436 691 449
rect 641 433 650 436
rect 617 432 641 433
rect 490 427 518 430
rect 1096 412 1099 415
rect 649 405 654 408
rect 712 404 744 407
rect 872 406 874 409
rect 487 393 490 401
rect 513 399 518 402
rect 639 399 654 402
rect 487 390 518 393
rect -3 314 0 317
rect -3 237 0 240
rect 487 188 490 390
rect 651 373 654 383
rect 688 380 691 388
rect 638 370 654 373
rect 498 283 501 294
rect 620 227 623 301
rect 706 258 712 261
rect 746 260 749 261
rect 671 255 674 256
rect 706 255 709 258
rect 695 252 709 255
rect 707 229 712 232
rect 770 228 776 231
rect 620 224 637 227
rect 695 223 712 226
rect 630 218 637 221
rect 613 199 616 210
rect 671 194 674 207
rect 692 202 695 207
rect 692 199 712 202
rect 746 199 749 212
rect 773 196 776 228
rect 1026 197 1029 200
rect 716 193 776 196
rect 487 185 496 188
rect 493 162 496 185
rect 575 183 579 186
rect 574 177 579 180
rect 637 178 640 181
rect 508 167 516 170
rect 574 169 577 177
rect 570 164 577 169
rect 713 167 719 170
rect 643 162 650 165
rect 643 152 646 162
rect 684 152 687 165
rect 713 152 716 167
rect 753 157 756 170
rect 637 149 646 152
rect 708 149 716 152
rect 613 148 637 149
rect 490 143 514 146
rect 799 138 805 141
rect 716 126 719 129
rect 799 128 802 138
rect 777 125 802 128
rect 645 121 650 124
rect 708 120 719 123
rect 487 109 490 117
rect 509 115 514 118
rect 635 115 650 118
rect 487 106 514 109
rect 647 89 650 99
rect 684 96 687 104
rect 705 101 719 104
rect 753 101 756 109
rect 634 86 650 89
rect -2 30 1 33
rect -2 -8 40 -5
rect 45 -8 828 -5
<< m2contact >>
rect 490 962 495 967
rect 500 732 505 737
rect 633 741 638 746
rect 633 686 638 691
rect 479 680 484 685
rect 496 680 501 685
rect 503 451 508 456
rect 644 460 649 465
rect 644 405 649 410
rect 508 399 513 404
rect 619 301 624 306
rect 497 294 502 299
rect 497 278 502 283
rect 625 216 630 221
rect 711 191 716 196
rect 503 167 508 172
rect 640 176 645 181
rect 492 157 497 162
rect 711 126 716 131
rect 640 121 645 126
rect 504 115 509 120
<< metal2 >>
rect 267 1199 296 1202
rect 267 1041 270 1199
rect 295 1120 298 1148
rect 295 1117 373 1120
rect 267 1038 484 1041
rect 481 1019 484 1038
rect 479 1014 484 1019
rect 481 979 484 987
rect 481 976 504 979
rect 479 735 484 738
rect 491 728 494 962
rect 501 737 504 976
rect 567 729 623 732
rect 491 725 499 728
rect 12 718 17 721
rect 480 694 483 706
rect 480 691 492 694
rect 480 599 483 680
rect 489 606 492 691
rect 496 685 499 725
rect 489 603 506 606
rect 480 596 499 599
rect 480 413 483 425
rect 496 420 499 596
rect 503 456 506 603
rect 496 417 511 420
rect 480 410 501 413
rect 498 299 501 410
rect 508 404 511 417
rect 620 306 623 729
rect 635 691 638 741
rect 646 410 649 460
rect 748 290 751 349
rect 480 287 751 290
rect 480 173 483 287
rect 498 272 501 278
rect 498 269 506 272
rect 503 172 506 269
rect 625 169 628 216
rect 574 166 628 169
rect 493 140 496 157
rect 493 137 508 140
rect 505 120 508 137
rect 642 126 645 176
rect 712 131 715 191
<< m123contact >>
rect 97 1270 102 1275
rect 546 1269 551 1274
rect 410 1261 415 1266
rect 257 1051 262 1056
rect 410 1143 415 1148
rect 373 1115 378 1120
rect 539 1036 544 1041
rect 612 993 617 998
rect 742 994 747 999
rect 537 970 542 975
rect 576 963 581 968
rect 549 773 554 778
rect 596 772 601 777
rect 563 748 568 753
rect 588 651 593 656
rect 597 651 602 656
rect 560 492 565 497
rect 609 489 614 494
rect 574 467 579 472
rect 599 370 604 375
rect 848 687 853 692
rect 628 677 633 682
rect 866 406 872 412
rect 665 253 670 258
rect 702 229 707 234
rect 1001 227 1006 232
rect 556 208 561 213
rect 613 194 618 199
rect 570 183 575 188
rect 805 191 810 196
rect 665 162 670 167
rect 595 86 600 91
rect 40 -9 45 -4
rect 828 -8 833 -3
<< metal3 >>
rect 98 1245 101 1270
rect 411 1148 414 1261
rect 547 1229 550 1269
rect 375 1053 378 1115
rect 411 1060 414 1143
rect 443 1067 446 1164
rect 501 1074 504 1112
rect 501 1071 832 1074
rect 443 1064 775 1067
rect 411 1057 746 1060
rect 258 1046 261 1051
rect 375 1050 705 1053
rect 258 1043 347 1046
rect 344 796 347 1043
rect 407 1043 542 1046
rect 407 1030 410 1043
rect 539 1041 542 1043
rect 539 966 542 970
rect 539 963 576 966
rect 539 937 542 963
rect 449 934 542 937
rect 344 793 567 796
rect 407 782 553 785
rect 407 749 410 782
rect 550 778 553 782
rect 564 753 567 793
rect 597 656 600 772
rect 449 653 588 656
rect 613 506 616 993
rect 407 501 564 504
rect 407 468 410 501
rect 561 497 564 501
rect 575 503 616 506
rect 575 472 578 503
rect 610 375 613 489
rect 449 372 599 375
rect 604 372 613 375
rect 629 334 632 677
rect 571 331 632 334
rect 407 217 560 220
rect 407 184 410 217
rect 557 213 560 217
rect 571 188 574 331
rect 449 91 450 92
rect 449 88 595 91
rect 614 89 617 194
rect 666 167 669 253
rect 702 234 705 1050
rect 743 999 746 1057
rect 743 755 746 994
rect 772 982 775 1064
rect 829 1034 832 1071
rect 772 806 775 958
rect 876 848 879 912
rect 876 845 939 848
rect 772 803 882 806
rect 743 752 852 755
rect 849 692 852 752
rect 757 544 760 648
rect 849 546 852 687
rect 879 674 882 803
rect 936 726 939 845
rect 982 547 985 604
rect 757 541 792 544
rect 849 543 870 546
rect 789 417 792 541
rect 867 412 870 543
rect 954 544 985 547
rect 954 445 957 544
rect 867 317 871 406
rect 805 314 871 317
rect 805 196 808 314
rect 898 306 901 369
rect 862 303 901 306
rect 862 171 865 303
rect 1002 232 1005 323
rect 600 86 617 89
rect 41 -4 44 46
rect 829 -3 832 154
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 292 0 1 1105
box -3 -9 349 129
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use nor  nor_0
timestamp 1618580541
transform 1 0 505 0 1 1000
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 539 0 1 993
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 572 0 1 999
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1618628987
transform 1 0 621 0 -1 1036
box -3 -9 349 129
use nand  nand_1
timestamp 1618580231
transform 1 0 572 0 -1 740
box 0 -35 34 27
use inv  inv_1
timestamp 1618579805
transform 1 0 606 0 -1 747
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 683
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 643 0 1 691
box 0 -30 34 39
use inv  inv_2
timestamp 1618579805
transform 1 0 677 0 1 684
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1618628987
transform 1 0 728 0 -1 728
box -3 -9 349 129
use nand  nand_2
timestamp 1618580231
transform 1 0 583 0 -1 459
box 0 -35 34 27
use inv  inv_3
timestamp 1618579805
transform 1 0 617 0 -1 466
box 0 -15 24 33
use cla  cla_1
timestamp 1618627066
transform 1 0 527 0 1 402
box -9 -46 112 95
use nor  nor_2
timestamp 1618580541
transform 1 0 654 0 1 410
box 0 -30 34 39
use inv  inv_4
timestamp 1618579805
transform 1 0 688 0 1 403
box 0 -15 24 33
use sumffo  sumffo_3
timestamp 1618628987
transform 1 0 747 0 -1 447
box -3 -9 349 129
use nand  nand_3
timestamp 1618580231
transform 1 0 579 0 -1 175
box 0 -35 34 27
use inv  inv_5
timestamp 1618579805
transform 1 0 613 0 -1 182
box 0 -15 24 33
use nand  nand_4
timestamp 1618580231
transform 1 0 637 0 1 229
box 0 -35 34 27
use inv  inv_7
timestamp 1618579805
transform 1 0 671 0 1 222
box 0 -15 24 33
use nand  nand_5
timestamp 1618580231
transform 1 0 712 0 1 234
box 0 -35 34 27
use inv  inv_8
timestamp 1618579805
transform 1 0 746 0 1 227
box 0 -15 24 33
use cla  cla_2
timestamp 1618627066
transform 1 0 523 0 1 118
box -9 -46 112 95
use nor  nor_3
timestamp 1618580541
transform 1 0 650 0 1 126
box 0 -30 34 39
use inv  inv_6
timestamp 1618579805
transform 1 0 684 0 1 119
box 0 -15 24 33
use nor  nor_4
timestamp 1618580541
transform 1 0 719 0 1 131
box 0 -30 34 39
use inv  inv_9
timestamp 1618579805
transform 1 0 753 0 1 124
box 0 -15 24 33
use ffo  ffo_0
timestamp 1618618535
transform 1 0 819 0 -1 199
box -14 -42 207 91
<< labels >>
rlabel metal1 -3 314 -3 317 3 y3in
rlabel metal1 -3 1153 -3 1156 3 cinin
rlabel metal1 -3 1083 -3 1086 3 x1in
rlabel metal1 -3 876 -3 879 3 y1in
rlabel metal1 -3 802 -3 805 3 x2in
rlabel metal1 -3 595 -3 598 3 y2in
rlabel metal1 -3 521 -3 524 3 x3in
rlabel metal1 -3 237 -3 240 3 x4in
rlabel metal1 -2 30 -2 33 3 y4in
rlabel metal1 -3 1252 -3 1255 3 clk
rlabel metal1 71 1271 71 1271 5 vdd!
rlabel metal1 19 -7 19 -7 1 gnd!
rlabel metal1 1080 693 1080 696 7 z3o
rlabel metal1 1099 412 1099 415 7 z4o
rlabel metal1 1029 197 1029 200 1 couto
rlabel metal1 644 1137 644 1140 7 z1o
rlabel metal1 971 1001 971 1004 7 z2o
<< end >>
