magic
tech scmos
timestamp 1618832345
<< metal1 >>
rect 0 1270 97 1273
rect 102 1270 525 1273
rect 3 1263 632 1266
rect 3 1256 6 1263
rect 241 1212 423 1215
rect 420 1165 423 1212
rect 420 1162 514 1165
rect 639 1160 643 1163
rect 490 989 498 992
rect 490 963 491 966
rect 518 732 519 735
rect 490 708 519 711
rect 487 674 490 682
rect 518 680 519 683
rect 487 671 519 674
<< m2contact >>
rect 498 987 503 992
rect 491 961 496 966
rect 513 732 518 737
rect 513 680 518 685
<< metal2 >>
rect 478 1216 518 1219
rect 478 1019 481 1216
rect 492 683 495 961
rect 500 735 503 987
rect 500 732 513 735
rect 492 680 513 683
<< m123contact >>
rect 97 1270 102 1275
rect 525 1270 530 1275
rect 632 1261 637 1266
rect 634 1160 639 1165
<< metal3 >>
rect 98 1245 101 1270
rect 526 1251 529 1270
rect 634 1165 637 1261
use ffipgarr  ffipgarr_0
timestamp 1618827105
transform 1 0 19 0 1 846
box -19 -846 471 410
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 517 0 1 1122
box -3 -9 349 129
use cla  cla_0
timestamp 1618627066
transform 1 0 528 0 1 683
box -9 -46 112 95
use cla  cla_1
timestamp 1618627066
transform 1 0 537 0 1 407
box -9 -46 112 95
use cla  cla_2
timestamp 1618627066
transform 1 0 527 0 1 121
box -9 -46 112 95
<< end >>
