* SPICE3 file created from cla.ext - technology: scmos

.option scale=0.09u

M1000 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=210 ps=144
M1001 vdd g1 n nand_0/w_0_0# pfet w=12 l=2
+  ad=420 pd=218 as=96 ps=40
M1002 n inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 n g1 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1005 inv_0/op inv_0/in vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1006 l p0 nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1007 nor_0/a_13_6# p1 vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 gnd p0 l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1009 l p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 inv_0/in g0 nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1011 nor_1/a_13_6# p1 vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 gnd g0 inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1013 inv_0/in p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd nor_0/w_0_0# 0.31fF
C1 g0 inv_0/in 0.16fF
C2 g1 inv_0/op 0.35fF
C3 n nand_0/w_0_0# 0.04fF
C4 gnd inv_0/op 0.10fF
C5 p1 vdd 0.15fF
C6 vdd l 0.20fF
C7 p1 g0 0.24fF
C8 vdd g1 0.07fF
C9 vdd gnd 0.33fF
C10 nor_1/w_0_0# vdd 0.31fF
C11 p1 inv_0/in 0.02fF
C12 n g1 0.13fF
C13 g0 g1 0.06fF
C14 gnd n 0.03fF
C15 vdd p0 0.06fF
C16 p1 nor_0/w_0_0# 0.06fF
C17 nor_1/w_0_0# g0 0.06fF
C18 inv_0/w_0_6# inv_0/op 0.03fF
C19 inv_0/in g1 0.04fF
C20 vdd inv_0/op 0.17fF
C21 l nor_0/w_0_0# 0.05fF
C22 inv_0/in gnd 0.30fF
C23 g1 nand_0/w_0_0# 0.06fF
C24 nor_1/w_0_0# inv_0/in 0.05fF
C25 p1 l 0.02fF
C26 inv_0/in inv_0/op 0.04fF
C27 p1 g1 0.00fF
C28 p0 nor_0/w_0_0# 0.06fF
C29 vdd inv_0/w_0_6# 0.06fF
C30 p1 gnd 0.50fF
C31 inv_0/op nand_0/w_0_0# 0.06fF
C32 p1 nor_1/w_0_0# 0.06fF
C33 l gnd 0.18fF
C34 vdd n 0.28fF
C35 vdd g0 0.06fF
C36 p1 p0 0.24fF
C37 gnd g1 0.20fF
C38 nor_1/w_0_0# g1 0.02fF
C39 l p0 0.16fF
C40 inv_0/in inv_0/w_0_6# 0.06fF
C41 vdd inv_0/in 0.05fF
C42 vdd nand_0/w_0_0# 0.10fF
C43 g0 Gnd 0.23fF
C44 p1 Gnd 0.53fF
C45 nor_1/w_0_0# Gnd 1.23fF
C46 l Gnd 0.06fF
C47 vdd Gnd 0.90fF
C48 p0 Gnd 0.18fF
C49 nor_0/w_0_0# Gnd 1.23fF
C50 inv_0/in Gnd 0.27fF
C51 inv_0/w_0_6# Gnd 0.58fF
C52 gnd Gnd 1.40fF
C53 n Gnd 0.09fF
C54 g1 Gnd 0.33fF
C55 inv_0/op Gnd 0.26fF
C56 nand_0/w_0_0# Gnd 0.82fF
