* SPICE3 file created from tspc.ext - technology: scmos

.option scale=0.01u

M1000 clk clk gnd Gnd nfet w=54 l=18
+  ad=2430 pd=198 as=17010 ps=1116
M1001 clk clk vdd inv_0/w_0_6# pfet w=108 l=18
+  ad=4860 pd=306 as=21870 ps=1332
M1002 a_n69_1# d gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1003 d a_13_35# vdd w_0_29# pfet w=126 l=18
+  ad=34020 pd=1044 as=0 ps=0
M1004 a_13_1# d gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1005 d clk a_n35_1# Gnd nfet w=108 l=18
+  ad=13608 pd=684 as=5832 ps=324
M1006 a_13_35# d vdd w_0_29# pfet w=126 l=18
+  ad=17010 pd=522 as=0 ps=0
M1007 a_13_35# clk a_13_1# Gnd nfet w=108 l=18
+  ad=6804 pd=342 as=0 ps=0
M1008 a_n35_1# a_n69_35# gnd Gnd nfet w=108 l=18
+  ad=0 pd=0 as=0 ps=0
M1009 a_n69_35# d vdd w_n82_29# pfet w=126 l=18
+  ad=17010 pd=522 as=0 ps=0
M1010 a_47_1# a_13_35# gnd Gnd nfet w=108 l=18
+  ad=5832 pd=324 as=0 ps=0
M1011 a_n69_35# clk a_n69_1# Gnd nfet w=108 l=18
+  ad=6804 pd=342 as=0 ps=0
M1012 d clk a_47_1# Gnd nfet w=108 l=18
+  ad=0 pd=0 as=0 ps=0
M1013 d a_n69_35# vdd w_n82_29# pfet w=126 l=18
+  ad=0 pd=0 as=0 ps=0
C0 a_n69_35# vdd 0.03fF
C1 clk d 0.98fF
C2 a_13_35# clk 0.46fF
C3 d vdd 0.13fF
C4 clk a_n69_1# 0.01fF
C5 a_13_35# vdd 0.03fF
C6 clk vdd 0.17fF
C7 a_n69_35# w_n82_29# 0.10fF
C8 d w_n82_29# 0.10fF
C9 a_n69_35# gnd 0.03fF
C10 d gnd 0.07fF
C11 a_13_35# gnd 0.03fF
C12 vdd w_n82_29# 0.14fF
C13 clk gnd 0.47fF
C14 inv_0/w_0_6# d 0.13fF
C15 w_0_29# d 0.10fF
C16 a_n35_1# clk 0.01fF
C17 w_0_29# a_13_35# 0.10fF
C18 clk inv_0/w_0_6# 0.31fF
C19 inv_0/w_0_6# vdd 0.06fF
C20 w_0_29# vdd 0.14fF
C21 a_n69_35# clk 0.54fF
C22 d Gnd 0.89fF
C23 w_0_29# Gnd 0.39fF
C24 w_n82_29# Gnd 0.39fF
C25 gnd Gnd 0.29fF
C26 clk Gnd 2.64fF
C27 vdd Gnd 0.18fF
C28 inv_0/w_0_6# Gnd 0.58fF
