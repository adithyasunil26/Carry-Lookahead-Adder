* SPICE3 file created from ffipgarrcla.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=11070 ps=6708
M1001 vdd nand_5/a inv_1/in inv_1/w_0_6# pfet w=12 l=2
+  ad=22140 pd=12236 as=96 ps=40
M1002 inv_1/in cla_0/l vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_1/in nand_5/a nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_2/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_0/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_2/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# nand_5/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd inv_7/op inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in nand_5/a vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in inv_7/op nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_0/g0 ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_0/g0 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1059 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1060 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1061 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1062 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1063 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1064 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_0/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op sumffo_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/ffi_1/q vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 nor_0/a ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1069 ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_0/ffi_0/q vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 gnd ffipgarr_0/ffipg_0/ffi_1/q nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1071 nor_0/a ffipgarr_0/ffipg_0/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1073 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1074 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1076 ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1077 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1078 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 ffipgarr_0/ffipg_0/ffi_0/nand_1/a clk ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# y1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1081 vdd clk ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1082 ffipgarr_0/ffipg_0/ffi_0/nand_3/a y1in vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 ffipgarr_0/ffipg_0/ffi_0/nand_3/a clk ffipgarr_0/ffipg_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1084 ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1085 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1086 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b ffipgarr_0/ffipg_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1088 ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1089 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1090 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1093 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1094 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 ffipgarr_0/ffipg_0/ffi_0/nand_7/a ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1096 ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1097 vdd ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1098 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1100 ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1101 vdd ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1102 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 ffipgarr_0/ffipg_0/ffi_0/inv_0/op y1in vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1107 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1108 ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1109 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1110 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1112 ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1113 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1114 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 ffipgarr_0/ffipg_0/ffi_1/nand_1/a clk ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1117 vdd clk ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1118 ffipgarr_0/ffipg_0/ffi_1/nand_3/a x1in vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 ffipgarr_0/ffipg_0/ffi_1/nand_3/a clk ffipgarr_0/ffipg_0/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1121 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1122 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1124 ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1125 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1126 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1128 ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1129 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1130 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1133 vdd ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1134 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1136 ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_0/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1137 vdd ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1138 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1140 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1141 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1142 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1145 vdd ffipgarr_0/ffipg_1/ffi_0/q cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1146 cla_1/g0 ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1148 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1153 sumffo_1/k ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1154 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1155 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1156 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_1/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op sumffo_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/ffi_1/q vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 cla_1/p0 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1161 ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_1/ffi_0/q vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 gnd ffipgarr_0/ffipg_1/ffi_1/q cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1163 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1165 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1166 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1168 ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1169 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1170 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ffipgarr_0/ffipg_1/ffi_0/nand_1/a clk ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1172 ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# y2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1173 vdd clk ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1174 ffipgarr_0/ffipg_1/ffi_0/nand_3/a y2in vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 ffipgarr_0/ffipg_1/ffi_0/nand_3/a clk ffipgarr_0/ffipg_1/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1176 ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1177 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1178 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1181 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1182 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1184 ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1185 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1186 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b ffipgarr_0/ffipg_1/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1188 ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1189 vdd ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1190 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1192 ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1193 vdd ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1194 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar ffipgarr_0/ffipg_1/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1196 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1197 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1201 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1202 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1204 ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1205 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1206 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipgarr_0/ffipg_1/ffi_1/nand_1/a clk ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1208 ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1209 vdd clk ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1210 ffipgarr_0/ffipg_1/ffi_1/nand_3/a x2in vdd ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 ffipgarr_0/ffipg_1/ffi_1/nand_3/a clk ffipgarr_0/ffipg_1/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1212 ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1213 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1214 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b ffipgarr_0/ffipg_1/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1216 ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1217 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1218 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1221 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1222 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1224 ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1225 vdd ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1226 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1228 ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_1/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1229 vdd ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1230 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1232 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1233 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1234 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1235 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1236 ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1237 vdd ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1238 cla_2/g0 ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 cla_2/g0 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1240 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1241 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1242 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1243 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1244 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1245 sumffo_2/k ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1246 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1247 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1248 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_2/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op sumffo_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_1/q vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1253 ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_2/ffi_0/q vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 gnd ffipgarr_0/ffipg_2/ffi_1/q cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1255 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1257 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1258 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1260 ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1261 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1262 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 ffipgarr_0/ffipg_2/ffi_0/nand_1/a clk ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1264 ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# y3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1265 vdd clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1266 ffipgarr_0/ffipg_2/ffi_0/nand_3/a y3in vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 ffipgarr_0/ffipg_2/ffi_0/nand_3/a clk ffipgarr_0/ffipg_2/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1268 ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1269 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1270 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1272 ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1273 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1274 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1276 ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1277 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1278 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1280 ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1281 vdd ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1282 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1284 ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1285 vdd ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1286 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar ffipgarr_0/ffipg_2/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1288 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1289 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1290 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1291 ffipgarr_0/ffipg_2/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1292 ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1293 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1294 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1296 ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1297 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1298 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 ffipgarr_0/ffipg_2/ffi_1/nand_1/a clk ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1300 ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1301 vdd clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1302 ffipgarr_0/ffipg_2/ffi_1/nand_3/a x3in vdd ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 ffipgarr_0/ffipg_2/ffi_1/nand_3/a clk ffipgarr_0/ffipg_2/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1304 ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1305 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1306 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1308 ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1309 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1310 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1312 ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1313 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1314 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b ffipgarr_0/ffipg_2/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1316 ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1317 vdd ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1318 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1320 ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_2/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1321 vdd ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1322 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar ffipgarr_0/ffipg_2/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1324 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1325 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1326 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1327 ffipgarr_0/ffipg_2/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1328 ffipgarr_0/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1329 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1330 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/a vdd ffipgarr_0/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1332 ffipgarr_0/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1333 vdd clk ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1334 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/inv_0/op vdd ffipgarr_0/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 ffipgarr_0/ffi_0/nand_1/a clk ffipgarr_0/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1336 ffipgarr_0/ffi_0/nand_2/a_13_n26# cinin gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1337 vdd clk ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1338 ffipgarr_0/ffi_0/nand_3/a cinin vdd ffipgarr_0/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 ffipgarr_0/ffi_0/nand_3/a clk ffipgarr_0/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1340 ffipgarr_0/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1341 vdd ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1342 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/a vdd ffipgarr_0/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1344 ffipgarr_0/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1345 vdd ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1346 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/nand_3/b vdd ffipgarr_0/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 ffipgarr_0/ffi_0/nand_6/a ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1348 ffipgarr_0/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1349 vdd ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1350 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/inv_1/op vdd ffipgarr_0/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1352 ffipgarr_0/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1353 vdd nand_5/a nor_0/b ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1354 nor_0/b ffipgarr_0/ffi_0/nand_6/a vdd ffipgarr_0/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 nor_0/b nand_5/a ffipgarr_0/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1356 ffipgarr_0/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1357 vdd nor_0/b nand_5/a ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1358 nand_5/a ffipgarr_0/ffi_0/nand_7/a vdd ffipgarr_0/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 nand_5/a nor_0/b ffipgarr_0/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1360 ffipgarr_0/ffi_0/inv_0/op cinin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1361 ffipgarr_0/ffi_0/inv_0/op cinin vdd ffipgarr_0/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1362 ffipgarr_0/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1363 ffipgarr_0/ffi_0/inv_1/op clk vdd ffipgarr_0/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1364 ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1365 vdd ffipgarr_0/ffipg_3/ffi_0/q cla_2/g1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1366 cla_2/g1 ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1368 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1369 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1370 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1371 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1372 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1373 sumffo_3/k ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1374 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1375 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1376 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_n43# ffipgarr_0/ffipg_3/ffi_1/q gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_38_n43# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_1/q vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1381 ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# ffipgarr_0/ffipg_3/ffi_0/q vdd ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 gnd ffipgarr_0/ffipg_3/ffi_1/q cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1383 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1385 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1386 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1388 ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1389 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1390 ffipgarr_0/ffipg_3/ffi_0/nand_1/a ffipgarr_0/ffipg_3/ffi_0/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ffipgarr_0/ffipg_3/ffi_0/nand_1/a clk ffipgarr_0/ffipg_3/ffi_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1392 ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# y4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1393 vdd clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1394 ffipgarr_0/ffipg_3/ffi_0/nand_3/a y4in vdd ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 ffipgarr_0/ffipg_3/ffi_0/nand_3/a clk ffipgarr_0/ffipg_3/ffi_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1396 ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1397 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1398 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1400 ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1401 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1402 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1404 ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1405 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1406 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1408 ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1409 vdd ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1410 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1412 ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1413 vdd ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1414 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1415 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1416 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1417 ffipgarr_0/ffipg_3/ffi_0/inv_0/op y4in vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1418 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1419 ffipgarr_0/ffipg_3/ffi_0/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1420 ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1421 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1422 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1424 ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1425 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1426 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/inv_0/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1427 ffipgarr_0/ffipg_3/ffi_1/nand_1/a clk ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1428 ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1429 vdd clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1430 ffipgarr_0/ffipg_3/ffi_1/nand_3/a x4in vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 ffipgarr_0/ffipg_3/ffi_1/nand_3/a clk ffipgarr_0/ffipg_3/ffi_1/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1432 ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1433 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1434 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1435 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1436 ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1437 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1438 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1440 ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/inv_1/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1441 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1442 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op vdd ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1443 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1444 ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1445 vdd ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1446 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1448 ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# ffipgarr_0/ffipg_3/ffi_1/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1449 vdd ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1450 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1451 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1452 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1453 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1454 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1455 ffipgarr_0/ffipg_3/ffi_1/inv_1/op clk vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1456 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1457 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1458 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1459 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1460 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1461 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1462 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1463 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1465 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1467 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1469 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1470 sumffo_0/ffo_0/nand_1/a_13_n26# sumffo_0/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1471 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1472 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/a vdd sumffo_0/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1474 sumffo_0/ffo_0/nand_0/a_13_n26# sumffo_0/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1475 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1476 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/inv_0/op vdd sumffo_0/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1478 sumffo_0/ffo_0/nand_2/a_13_n26# sumffo_0/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1479 vdd sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1480 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 sumffo_0/ffo_0/nand_3/a sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1482 sumffo_0/ffo_0/nand_3/a_13_n26# sumffo_0/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1483 vdd sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1484 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/a vdd sumffo_0/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1486 sumffo_0/ffo_0/nand_4/a_13_n26# sumffo_0/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1487 vdd clk sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1488 sumffo_0/ffo_0/nand_6/a sumffo_0/ffo_0/nand_3/b vdd sumffo_0/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 sumffo_0/ffo_0/nand_6/a clk sumffo_0/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1490 sumffo_0/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1491 vdd sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1492 sumffo_0/ffo_0/nand_7/a clk vdd sumffo_0/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1494 sumffo_0/ffo_0/nand_6/a_13_n26# sumffo_0/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1495 vdd z1o sumffo_0/sbar sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1496 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a vdd sumffo_0/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 sumffo_0/sbar z1o sumffo_0/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1498 sumffo_0/ffo_0/nand_7/a_13_n26# sumffo_0/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1499 vdd sumffo_0/sbar z1o sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1500 z1o sumffo_0/ffo_0/nand_7/a vdd sumffo_0/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 z1o sumffo_0/sbar sumffo_0/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1502 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1503 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d vdd sumffo_0/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1504 sumffo_0/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1505 sumffo_0/ffo_0/nand_0/b clk vdd sumffo_0/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1506 sumffo_0/xor_0/inv_0/op sumffo_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1507 sumffo_0/xor_0/inv_0/op sumffo_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1508 sumffo_0/xor_0/inv_1/op nand_5/a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1509 sumffo_0/xor_0/inv_1/op nand_5/a vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1510 vdd nand_5/a sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1511 sumffo_0/ffo_0/d nand_5/a sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1512 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1513 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op sumffo_0/ffo_0/d sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1514 sumffo_0/xor_0/a_10_n43# sumffo_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1515 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op sumffo_0/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 sumffo_0/xor_0/a_10_10# sumffo_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 sumffo_2/ffo_0/nand_1/a_13_n26# sumffo_2/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1519 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1520 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a vdd sumffo_2/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1521 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1522 sumffo_2/ffo_0/nand_0/a_13_n26# sumffo_2/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1523 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1524 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/inv_0/op vdd sumffo_2/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1526 sumffo_2/ffo_0/nand_2/a_13_n26# sumffo_2/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1527 vdd sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1528 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1529 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1530 sumffo_2/ffo_0/nand_3/a_13_n26# sumffo_2/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1531 vdd sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1532 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/a vdd sumffo_2/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1534 sumffo_2/ffo_0/nand_4/a_13_n26# sumffo_2/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1535 vdd clk sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1536 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_3/b vdd sumffo_2/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 sumffo_2/ffo_0/nand_6/a clk sumffo_2/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1538 sumffo_2/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1539 vdd sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1540 sumffo_2/ffo_0/nand_7/a clk vdd sumffo_2/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1541 sumffo_2/ffo_0/nand_7/a sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1542 sumffo_2/ffo_0/nand_6/a_13_n26# sumffo_2/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1543 vdd z3o sumffo_2/sbar sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1544 sumffo_2/sbar sumffo_2/ffo_0/nand_6/a vdd sumffo_2/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 sumffo_2/sbar z3o sumffo_2/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1546 sumffo_2/ffo_0/nand_7/a_13_n26# sumffo_2/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1547 vdd sumffo_2/sbar z3o sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1548 z3o sumffo_2/ffo_0/nand_7/a vdd sumffo_2/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 z3o sumffo_2/sbar sumffo_2/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1550 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1551 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d vdd sumffo_2/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1552 sumffo_2/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1553 sumffo_2/ffo_0/nand_0/b clk vdd sumffo_2/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1554 sumffo_2/xor_0/inv_0/op sumffo_2/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1555 sumffo_2/xor_0/inv_0/op sumffo_2/k vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1556 sumffo_2/xor_0/inv_1/op inv_2/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1557 sumffo_2/xor_0/inv_1/op inv_2/op vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1558 vdd inv_2/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1559 sumffo_2/ffo_0/d inv_2/op sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1560 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1561 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1562 sumffo_2/xor_0/a_10_n43# sumffo_2/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 sumffo_2/xor_0/a_10_10# sumffo_2/k vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1565 sumffo_2/ffo_0/d sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 sumffo_1/ffo_0/nand_1/a_13_n26# sumffo_1/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1567 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1568 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a vdd sumffo_1/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1570 sumffo_1/ffo_0/nand_0/a_13_n26# sumffo_1/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1571 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1572 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/inv_0/op vdd sumffo_1/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1573 sumffo_1/ffo_0/nand_1/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1574 sumffo_1/ffo_0/nand_2/a_13_n26# sumffo_1/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1575 vdd sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1576 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1578 sumffo_1/ffo_0/nand_3/a_13_n26# sumffo_1/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1579 vdd sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1580 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/a vdd sumffo_1/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1582 sumffo_1/ffo_0/nand_4/a_13_n26# sumffo_1/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1583 vdd clk sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1584 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_3/b vdd sumffo_1/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1585 sumffo_1/ffo_0/nand_6/a clk sumffo_1/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1586 sumffo_1/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1587 vdd sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1588 sumffo_1/ffo_0/nand_7/a clk vdd sumffo_1/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1590 sumffo_1/ffo_0/nand_6/a_13_n26# sumffo_1/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1591 vdd z2o sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1592 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a vdd sumffo_1/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 sumffo_1/sbar z2o sumffo_1/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1594 sumffo_1/ffo_0/nand_7/a_13_n26# sumffo_1/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1595 vdd sumffo_1/sbar z2o sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1596 z2o sumffo_1/ffo_0/nand_7/a vdd sumffo_1/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 z2o sumffo_1/sbar sumffo_1/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1598 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1599 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d vdd sumffo_1/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1600 sumffo_1/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1601 sumffo_1/ffo_0/nand_0/b clk vdd sumffo_1/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1602 sumffo_1/xor_0/inv_0/op sumffo_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1603 sumffo_1/xor_0/inv_0/op sumffo_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1604 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1605 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1606 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1607 sumffo_1/ffo_0/d nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1608 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1609 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op sumffo_1/ffo_0/d sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1610 sumffo_1/xor_0/a_10_n43# sumffo_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1611 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 sumffo_1/xor_0/a_10_10# sumffo_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1614 sumffo_3/ffo_0/nand_1/a_13_n26# sumffo_3/ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1615 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1616 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/a vdd sumffo_3/ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1618 sumffo_3/ffo_0/nand_0/a_13_n26# sumffo_3/ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1619 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1620 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/inv_0/op vdd sumffo_3/ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1622 sumffo_3/ffo_0/nand_2/a_13_n26# sumffo_3/ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1623 vdd sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1624 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1626 sumffo_3/ffo_0/nand_3/a_13_n26# sumffo_3/ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1627 vdd sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1628 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/a vdd sumffo_3/ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1630 sumffo_3/ffo_0/nand_4/a_13_n26# sumffo_3/ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1631 vdd clk sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1632 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_3/b vdd sumffo_3/ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 sumffo_3/ffo_0/nand_6/a clk sumffo_3/ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1634 sumffo_3/ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1635 vdd sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1636 sumffo_3/ffo_0/nand_7/a clk vdd sumffo_3/ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 sumffo_3/ffo_0/nand_7/a sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1638 sumffo_3/ffo_0/nand_6/a_13_n26# sumffo_3/ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1639 vdd z4o sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1640 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a vdd sumffo_3/ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 sumffo_3/sbar z4o sumffo_3/ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1642 sumffo_3/ffo_0/nand_7/a_13_n26# sumffo_3/ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1643 vdd sumffo_3/sbar z4o sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1644 z4o sumffo_3/ffo_0/nand_7/a vdd sumffo_3/ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1645 z4o sumffo_3/sbar sumffo_3/ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1646 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1647 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/d vdd sumffo_3/ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1648 sumffo_3/ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1649 sumffo_3/ffo_0/nand_0/b clk vdd sumffo_3/ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1650 sumffo_3/xor_0/inv_0/op sumffo_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1651 sumffo_3/xor_0/inv_0/op sumffo_3/k vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1652 sumffo_3/xor_0/inv_1/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1653 sumffo_3/xor_0/inv_1/op inv_4/op vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1654 vdd inv_4/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1655 sumffo_3/ffo_0/d inv_4/op sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1656 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1657 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1658 sumffo_3/xor_0/a_10_n43# sumffo_3/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op sumffo_3/ffo_0/d Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 sumffo_3/xor_0/a_10_10# sumffo_3/k vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1662 ffo_0/nand_1/a_13_n26# ffo_0/nand_1/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1663 vdd ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1664 ffo_0/nand_3/b ffo_0/nand_1/a vdd ffo_0/nand_1/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1665 ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1666 ffo_0/nand_0/a_13_n26# ffo_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1667 vdd ffo_0/nand_0/b ffo_0/nand_1/a ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1668 ffo_0/nand_1/a ffo_0/inv_0/op vdd ffo_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 ffo_0/nand_1/a ffo_0/nand_0/b ffo_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1670 ffo_0/nand_2/a_13_n26# ffo_0/d gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1671 vdd ffo_0/nand_0/b ffo_0/nand_3/a ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1672 ffo_0/nand_3/a ffo_0/d vdd ffo_0/nand_2/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1673 ffo_0/nand_3/a ffo_0/nand_0/b ffo_0/nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1674 ffo_0/nand_3/a_13_n26# ffo_0/nand_3/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1675 vdd ffo_0/nand_3/b ffo_0/nand_1/b ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1676 ffo_0/nand_1/b ffo_0/nand_3/a vdd ffo_0/nand_3/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 ffo_0/nand_1/b ffo_0/nand_3/b ffo_0/nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1678 ffo_0/nand_4/a_13_n26# ffo_0/nand_3/b gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1679 vdd clk ffo_0/nand_6/a ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1680 ffo_0/nand_6/a ffo_0/nand_3/b vdd ffo_0/nand_4/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ffo_0/nand_6/a clk ffo_0/nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1682 ffo_0/nand_5/a_13_n26# clk gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1683 vdd ffo_0/nand_1/b ffo_0/nand_7/a ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1684 ffo_0/nand_7/a clk vdd ffo_0/nand_5/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ffo_0/nand_7/a ffo_0/nand_1/b ffo_0/nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1686 ffo_0/nand_6/a_13_n26# ffo_0/nand_6/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1687 vdd couto ffo_0/qbar ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1688 ffo_0/qbar ffo_0/nand_6/a vdd ffo_0/nand_6/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 ffo_0/qbar couto ffo_0/nand_6/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1690 ffo_0/nand_7/a_13_n26# ffo_0/nand_7/a gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1691 vdd ffo_0/qbar couto ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1692 couto ffo_0/nand_7/a vdd ffo_0/nand_7/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1693 couto ffo_0/qbar ffo_0/nand_7/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1694 ffo_0/inv_0/op ffo_0/d gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1695 ffo_0/inv_0/op ffo_0/d vdd ffo_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1696 ffo_0/nand_0/b clk gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1697 ffo_0/nand_0/b clk vdd ffo_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1698 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1699 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1700 nor_1/b inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1701 nor_1/b inv_1/in vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1702 inv_2/op inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1703 inv_2/op inv_2/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1704 inv_0/in nor_0/b nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1705 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1706 gnd nor_0/b inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1707 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1708 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1709 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1710 inv_2/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1711 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 gnd nor_1/b inv_2/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1713 inv_2/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1714 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1715 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1716 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1717 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1719 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 nor_4/a inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1721 nor_4/a inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1722 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1723 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1724 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1725 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1726 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1727 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1728 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1729 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1730 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1731 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1732 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1733 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1734 nor_4/b inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1735 nor_4/b inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1736 ffo_0/d inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1737 ffo_0/d inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
C0 ffipgarr_0/ffipg_0/ffi_1/inv_1/op x1in 0.01fF
C1 vdd cla_1/nor_0/a_13_6# 0.01fF
C2 vdd inv_0/in 0.09fF
C3 vdd ffo_0/nand_3/w_0_0# 0.11fF
C4 sumffo_1/xor_0/inv_1/w_0_6# nand_2/b 0.23fF
C5 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C6 z2o sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C7 vdd sumffo_0/ffo_0/nand_4/w_0_0# 0.10fF
C8 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C9 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C10 cla_0/inv_0/w_0_6# cla_0/inv_0/in 0.06fF
C11 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/w_0_0# 0.04fF
C12 sumffo_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C13 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/b 0.32fF
C14 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/op 1.63fF
C15 vdd ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.10fF
C16 vdd inv_3/in 0.30fF
C17 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_1/a 0.04fF
C18 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C19 ffo_0/nand_7/a gnd 0.03fF
C20 vdd cla_2/p1 0.31fF
C21 cla_1/p0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C22 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# y1in 0.06fF
C23 ffo_0/nand_3/a ffo_0/nand_3/b 0.31fF
C24 sumffo_3/ffo_0/nand_6/w_0_0# sumffo_3/ffo_0/nand_6/a 0.06fF
C25 clk sumffo_2/ffo_0/nand_0/b 0.04fF
C26 gnd sumffo_2/ffo_0/inv_0/op 0.10fF
C27 ffipgarr_0/ffipg_3/ffi_0/nand_7/a ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.06fF
C28 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.04fF
C29 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.31fF
C30 ffo_0/d ffo_0/nand_2/w_0_0# 0.06fF
C31 sumffo_1/k sumffo_1/xor_0/w_n3_4# 0.06fF
C32 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C33 sumffo_2/ffo_0/inv_1/w_0_6# clk 0.06fF
C34 vdd sumffo_2/sbar 0.28fF
C35 vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.10fF
C36 vdd ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C37 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.21fF
C38 ffo_0/nand_4/w_0_0# clk 0.06fF
C39 gnd inv_2/in 0.24fF
C40 cla_0/g0 gnd 0.94fF
C41 cla_2/p0 sumffo_3/k 0.09fF
C42 vdd z2o 0.28fF
C43 sumffo_2/k sumffo_2/xor_0/inv_0/w_0_6# 0.06fF
C44 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C45 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.15fF
C46 vdd nand_0/w_0_0# 0.10fF
C47 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/sbar 0.06fF
C48 vdd inv_1/in 0.30fF
C49 nor_3/b cla_2/l 0.27fF
C50 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C51 gnd ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.10fF
C52 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.31fF
C53 vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.10fF
C54 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_3/a 0.04fF
C55 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_6/w_0_0# 0.06fF
C56 gnd ffo_0/nand_1/a 0.03fF
C57 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C58 gnd sumffo_2/ffo_0/nand_1/a_13_n26# 0.01fF
C59 cla_0/nand_0/w_0_0# gnd 0.01fF
C60 ffipgarr_0/ffi_0/nand_6/w_0_0# nand_5/a 0.06fF
C61 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.04fF
C62 ffo_0/d ffo_0/nand_0/b 0.40fF
C63 sumffo_2/ffo_0/nand_6/a z3o 0.31fF
C64 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.00fF
C65 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# clk 0.06fF
C66 vdd x1in 0.04fF
C67 gnd ffipgarr_0/ffipg_2/ffi_0/nand_0/a_13_n26# 0.01fF
C68 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# gnd 0.00fF
C69 sumffo_2/ffo_0/nand_3/b gnd 0.52fF
C70 ffo_0/nand_0/w_0_0# ffo_0/inv_0/op 0.06fF
C71 gnd ffo_0/nand_3/b 0.35fF
C72 y4in ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C73 nor_0/b ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C74 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.06fF
C75 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.06fF
C76 gnd ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.15fF
C77 nor_4/b nor_4/w_0_0# 0.06fF
C78 ffo_0/nand_7/a ffo_0/qbar 0.31fF
C79 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_0/op 0.06fF
C80 ffipgarr_0/ffi_0/inv_1/w_0_6# ffipgarr_0/ffi_0/inv_1/op 0.04fF
C81 cla_2/p0 ffipgarr_0/ffipg_2/ffi_0/q 0.03fF
C82 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.04fF
C83 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C84 sumffo_2/ffo_0/nand_0/w_0_0# cla_0/n 0.04fF
C85 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_1/a 0.13fF
C86 vdd sumffo_1/ffo_0/nand_6/a 0.30fF
C87 vdd sumffo_2/ffo_0/nand_7/a 0.30fF
C88 cla_2/g0 cla_1/n 0.13fF
C89 gnd ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.22fF
C90 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/qbar 0.31fF
C91 gnd ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.03fF
C92 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/inv_0/op 0.03fF
C93 vdd ffipgarr_0/ffipg_3/ffi_0/qbar 0.33fF
C94 ffipgarr_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.04fF
C95 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C96 vdd ffipgarr_0/ffipg_1/ffi_0/q 0.38fF
C97 ffipgarr_0/ffipg_0/ffi_0/inv_0/op clk 0.32fF
C98 cla_0/nor_1/w_0_0# cla_1/p0 0.06fF
C99 cla_0/nand_0/a_13_n26# nand_2/b 0.00fF
C100 sumffo_0/ffo_0/nand_6/w_0_0# z1o 0.06fF
C101 vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.34fF
C102 cla_0/l cla_2/g0 0.08fF
C103 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# gnd 0.00fF
C104 sumffo_1/ffo_0/nand_1/b sumffo_1/ffo_0/nand_1/a 0.31fF
C105 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.04fF
C106 cla_0/g0 nor_0/a 1.58fF
C107 ffo_0/inv_1/w_0_6# vdd 0.06fF
C108 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/b 0.32fF
C109 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.04fF
C110 vdd sumffo_3/xor_0/inv_0/w_0_6# 0.09fF
C111 vdd sumffo_0/xor_0/inv_1/w_0_6# 0.06fF
C112 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.04fF
C113 cla_2/nor_1/a_13_6# gnd 0.01fF
C114 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/w_0_0# 0.06fF
C115 vdd y4in 0.04fF
C116 vdd ffipgarr_0/ffi_0/nand_6/a 0.30fF
C117 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C118 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.27fF
C119 vdd ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.10fF
C120 vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.17fF
C121 vdd sumffo_2/ffo_0/nand_2/w_0_0# 0.10fF
C122 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/w_0_0# 0.06fF
C123 clk sumffo_0/ffo_0/nand_0/b 0.04fF
C124 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# clk 0.06fF
C125 cla_2/g1 gnd 0.27fF
C126 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.06fF
C127 gnd ffipgarr_0/ffipg_1/ffi_0/inv_1/op 0.22fF
C128 vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C129 cla_2/g1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C130 cinin ffipgarr_0/ffi_0/inv_1/op 0.01fF
C131 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.00fF
C132 y2in clk 0.70fF
C133 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C134 vdd sumffo_3/ffo_0/nand_6/a 0.30fF
C135 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/inv_0/op 0.32fF
C136 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C137 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/ffi_0/nand_0/w_0_0# 0.06fF
C138 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C139 clk cla_0/n 0.12fF
C140 sumffo_3/k inv_4/op 0.09fF
C141 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/a 0.00fF
C142 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.04fF
C143 cla_2/g0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C144 ffipgarr_0/ffipg_1/ffi_1/nand_3/a clk 0.13fF
C145 cla_1/p0 cla_1/l 0.16fF
C146 sumffo_3/xor_0/a_10_10# inv_4/op 0.12fF
C147 vdd inv_8/w_0_6# 0.15fF
C148 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C149 vdd x4in 0.04fF
C150 sumffo_1/k vdd 0.26fF
C151 vdd cla_0/inv_0/in 0.05fF
C152 gnd ffipgarr_0/ffipg_1/ffi_1/qbar 0.34fF
C153 inv_7/w_0_6# inv_7/in 0.10fF
C154 cla_0/nor_1/w_0_0# gnd 0.01fF
C155 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_1/op 0.52fF
C156 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.45fF
C157 gnd ffipgarr_0/ffi_0/inv_1/op 0.22fF
C158 ffipgarr_0/ffipg_2/ffi_1/nand_3/a ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.04fF
C159 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.06fF
C160 sumffo_3/xor_0/inv_1/w_0_6# inv_4/op 0.23fF
C161 vdd ffo_0/nand_1/b 0.31fF
C162 z1o sumffo_0/ffo_0/nand_7/w_0_0# 0.04fF
C163 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C164 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C165 vdd sumffo_3/ffo_0/nand_3/a 0.30fF
C166 x3in ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.01fF
C167 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C168 ffipgarr_0/ffipg_1/ffi_1/qbar ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C169 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.04fF
C170 ffipgarr_0/ffi_0/nand_2/w_0_0# cinin 0.06fF
C171 vdd ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# 0.10fF
C172 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# 0.45fF
C173 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# clk 0.06fF
C174 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C175 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C176 x4in ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C177 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.32fF
C178 vdd ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.17fF
C179 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.04fF
C180 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C181 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/w_n3_4# 0.06fF
C182 gnd sumffo_2/ffo_0/nand_1/b 0.38fF
C183 sumffo_0/ffo_0/inv_1/w_0_6# clk 0.06fF
C184 gnd ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.03fF
C185 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# 0.06fF
C186 cla_0/inv_0/op gnd 0.15fF
C187 sumffo_2/ffo_0/d sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C188 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.16fF
C189 vdd sumffo_3/ffo_0/nand_3/b 0.39fF
C190 ffo_0/nand_4/w_0_0# ffo_0/nand_3/b 0.06fF
C191 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_0/b 0.06fF
C192 sumffo_2/k sumffo_2/xor_0/w_n3_4# 0.06fF
C193 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C194 gnd ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.03fF
C195 cla_1/p0 gnd 0.74fF
C196 ffo_0/inv_0/w_0_6# gnd 0.01fF
C197 vdd ffo_0/nand_0/w_0_0# 0.10fF
C198 gnd sumffo_1/sbar 0.34fF
C199 vdd sumffo_1/ffo_0/nand_0/w_0_0# 0.10fF
C200 vdd ffipgarr_0/ffipg_1/ffi_0/qbar 0.33fF
C201 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.45fF
C202 cla_0/n sumffo_2/ffo_0/nand_1/a 0.08fF
C203 gnd sumffo_2/ffo_0/nand_1/w_0_0# 0.00fF
C204 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/nand_0/w_0_0# 0.06fF
C205 sumffo_1/xor_0/inv_0/op sumffo_1/ffo_0/d 0.06fF
C206 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_6/a 0.04fF
C207 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.04fF
C208 clk x3in 0.70fF
C209 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.06fF
C210 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.04fF
C211 vdd ffipgarr_0/ffipg_3/ffi_1/q 1.35fF
C212 clk y3in 0.70fF
C213 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.31fF
C214 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/a 0.30fF
C215 sumffo_1/ffo_0/d sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C216 gnd ffo_0/nand_3/a 0.14fF
C217 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.04fF
C218 gnd cla_1/l 0.18fF
C219 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.04fF
C220 gnd ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.14fF
C221 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.45fF
C222 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.75fF
C223 ffipgarr_0/ffipg_1/ffi_1/nand_7/a ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.06fF
C224 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.93fF
C225 inv_1/in nand_5/a 0.13fF
C226 clk sumffo_3/ffo_0/nand_1/b 0.45fF
C227 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# clk 0.06fF
C228 vdd ffipgarr_0/ffipg_3/ffi_0/q 0.38fF
C229 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C230 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C231 gnd sumffo_0/ffo_0/d 0.37fF
C232 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.33fF
C233 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C234 vdd ffipgarr_0/ffipg_2/ffi_1/qbar 0.33fF
C235 vdd ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# 0.10fF
C236 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C237 vdd cla_2/g0 0.45fF
C238 cla_0/l inv_7/w_0_6# 0.06fF
C239 gnd sumffo_1/ffo_0/nand_0/b 0.45fF
C240 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_3/w_0_0# 0.04fF
C241 y4in ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C242 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# vdd 0.10fF
C243 ffipgarr_0/ffipg_3/ffi_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.03fF
C244 ffipgarr_0/ffipg_0/ffi_1/inv_0/op clk 0.32fF
C245 sumffo_2/xor_0/inv_0/op inv_2/op 0.20fF
C246 gnd sumffo_0/ffo_0/nand_3/b 0.35fF
C247 gnd cinin 0.19fF
C248 gnd y1in 0.19fF
C249 sumffo_2/k cla_1/p0 2.09fF
C250 clk sumffo_0/ffo_0/nand_4/w_0_0# 0.06fF
C251 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C252 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.13fF
C253 sumffo_1/k sumffo_1/xor_0/inv_0/w_0_6# 0.06fF
C254 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_1/b 0.31fF
C255 vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.17fF
C256 clk ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.07fF
C257 ffipgarr_0/ffipg_2/ffi_0/nand_1/a ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C258 sumffo_0/k ffipgarr_0/ffipg_0/ffi_1/q 1.58fF
C259 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C260 gnd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.00fF
C261 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C262 ffipgarr_0/ffipg_1/ffi_0/nand_7/a gnd 0.03fF
C263 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.04fF
C264 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.13fF
C265 nor_3/b inv_6/in 0.16fF
C266 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_3/a 0.31fF
C267 sumffo_0/xor_0/w_n3_4# sumffo_0/k 0.06fF
C268 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/w_0_0# 0.04fF
C269 vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.17fF
C270 inv_1/w_0_6# cla_0/l 0.28fF
C271 sumffo_2/xor_0/inv_0/op vdd 0.15fF
C272 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.31fF
C273 gnd ffipgarr_0/ffipg_3/ffi_1/nand_0/a_13_n26# 0.01fF
C274 cla_0/n inv_2/in 0.02fF
C275 nor_1/b inv_1/w_0_6# 0.03fF
C276 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.04fF
C277 sumffo_3/sbar sumffo_3/ffo_0/nand_7/a 0.31fF
C278 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_1/op 0.08fF
C279 ffipgarr_0/ffipg_0/ffi_1/nand_7/a ffipgarr_0/ffipg_0/ffi_1/qbar 0.31fF
C280 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C281 cla_1/p0 nor_0/a 0.24fF
C282 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.06fF
C283 inv_8/w_0_6# nor_4/b 0.03fF
C284 ffo_0/nand_0/b ffo_0/inv_0/op 0.32fF
C285 vdd sumffo_1/ffo_0/nand_1/b 0.31fF
C286 nand_5/a sumffo_0/xor_0/inv_1/w_0_6# 0.23fF
C287 sumffo_0/ffo_0/d sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C288 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.31fF
C289 ffipgarr_0/ffi_0/nand_7/a nor_0/b 0.31fF
C290 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.39fF
C291 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C292 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.39fF
C293 z2o sumffo_1/ffo_0/nand_7/a 0.00fF
C294 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.04fF
C295 nand_5/a ffipgarr_0/ffi_0/nand_6/a 0.31fF
C296 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# gnd 0.00fF
C297 gnd ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.14fF
C298 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C299 x1in clk 0.70fF
C300 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C301 vdd inv_9/in 0.09fF
C302 vdd nor_0/b 0.90fF
C303 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C304 cla_2/inv_0/in cla_2/p1 0.02fF
C305 sumffo_2/k gnd 0.35fF
C306 nor_1/b nor_1/w_0_0# 0.06fF
C307 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.06fF
C308 sumffo_2/ffo_0/nand_3/b cla_0/n 0.19fF
C309 gnd sumffo_1/ffo_0/nand_0/a_13_n26# 0.01fF
C310 vdd sumffo_1/xor_0/inv_0/op 0.15fF
C311 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_3/a 0.13fF
C312 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C313 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.31fF
C314 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_1/q 0.27fF
C315 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.06fF
C316 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C317 clk sumffo_1/ffo_0/nand_6/a 0.13fF
C318 vdd sumffo_1/ffo_0/nand_2/w_0_0# 0.10fF
C319 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_4/w_0_0# 0.04fF
C320 vdd sumffo_0/xor_0/inv_0/w_0_6# 0.09fF
C321 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 1.63fF
C322 vdd ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.10fF
C323 ffo_0/qbar gnd 0.34fF
C324 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.04fF
C325 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C326 gnd ffipgarr_0/ffipg_0/ffi_0/qbar 0.34fF
C327 nand_5/a inv_8/w_0_6# 0.57fF
C328 sumffo_2/ffo_0/d sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C329 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/q 0.31fF
C330 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/ffi_0/q 0.20fF
C331 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.13fF
C332 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.04fF
C333 sumffo_1/k nand_5/a 0.02fF
C334 vdd sumffo_3/ffo_0/d 0.04fF
C335 vdd sumffo_1/ffo_0/nand_3/b 0.39fF
C336 z1o sumffo_0/ffo_0/nand_7/a 0.00fF
C337 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C338 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/inv_0/w_0_6# 0.03fF
C339 gnd ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.26fF
C340 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C341 ffo_0/inv_1/w_0_6# clk 0.06fF
C342 gnd ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.03fF
C343 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.04fF
C344 gnd nor_0/a 0.29fF
C345 cla_0/g0 cla_1/g0 0.18fF
C346 cla_0/l nand_2/b 0.46fF
C347 vdd sumffo_3/xor_0/inv_0/op 0.15fF
C348 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C349 nand_2/b sumffo_1/xor_0/w_n3_4# 0.06fF
C350 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.10fF
C351 vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C352 vdd cla_1/nor_1/w_0_0# 0.31fF
C353 ffipgarr_0/ffipg_2/ffi_0/inv_0/op y3in 0.04fF
C354 gnd sumffo_1/ffo_0/nand_3/a 0.03fF
C355 sumffo_3/sbar sumffo_3/ffo_0/nand_6/w_0_0# 0.04fF
C356 ffipgarr_0/ffipg_3/ffi_1/nand_7/a ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C357 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.06fF
C358 y4in clk 0.64fF
C359 ffipgarr_0/ffipg_1/ffi_0/inv_1/op y2in 0.01fF
C360 vdd sumffo_0/ffo_0/nand_1/a 0.30fF
C361 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C362 vdd inv_7/w_0_6# 0.20fF
C363 ffo_0/nand_6/w_0_0# ffo_0/nand_6/a 0.06fF
C364 clk ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.32fF
C365 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C366 sumffo_1/ffo_0/d sumffo_1/xor_0/inv_1/op 0.52fF
C367 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/a 0.06fF
C368 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.31fF
C369 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.39fF
C370 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C371 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C372 gnd ffipgarr_0/ffipg_2/ffi_1/q 0.93fF
C373 cla_2/l gnd 0.36fF
C374 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C375 clk sumffo_3/ffo_0/nand_6/a 0.13fF
C376 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C377 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# x2in 0.06fF
C378 cla_1/g0 cla_0/nand_0/w_0_0# 0.06fF
C379 vdd cla_0/nor_0/a_13_6# 0.01fF
C380 vdd ffo_0/nand_2/w_0_0# 0.10fF
C381 vdd sumffo_0/xor_0/inv_0/op 0.15fF
C382 vdd ffipgarr_0/ffi_0/nand_0/w_0_0# 0.10fF
C383 sumffo_3/sbar sumffo_3/ffo_0/nand_7/w_0_0# 0.06fF
C384 gnd sumffo_2/ffo_0/nand_0/b 0.38fF
C385 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C386 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C387 vdd nor_4/a 0.15fF
C388 ffo_0/nand_6/w_0_0# couto 0.06fF
C389 sumffo_3/ffo_0/nand_6/a z4o 0.31fF
C390 vdd sumffo_0/ffo_0/nand_3/a 0.30fF
C391 clk x4in 0.70fF
C392 vdd ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.11fF
C393 inv_1/w_0_6# vdd 0.15fF
C394 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# nand_5/a 0.04fF
C395 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/a_10_10# 0.16fF
C396 cla_1/inv_0/op gnd 0.15fF
C397 nand_0/w_0_0# cla_0/g0 0.06fF
C398 clk ffo_0/nand_1/b 0.45fF
C399 vdd ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C400 cla_1/g0 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C401 gnd ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.03fF
C402 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.12fF
C403 vdd inv_0/op 0.17fF
C404 inv_2/op nor_1/w_0_0# 0.03fF
C405 vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.34fF
C406 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/nand_5/w_0_0# 0.06fF
C407 sumffo_2/k ffipgarr_0/ffipg_2/ffi_1/q 2.17fF
C408 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C409 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C410 cla_0/l sumffo_3/k 0.06fF
C411 vdd sumffo_2/ffo_0/nand_6/w_0_0# 0.10fF
C412 gnd ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.35fF
C413 ffo_0/nand_3/b ffo_0/nand_3/w_0_0# 0.06fF
C414 vdd ffo_0/nand_0/b 0.15fF
C415 sumffo_2/xor_0/inv_1/w_0_6# inv_2/op 0.23fF
C416 z1o sumffo_0/sbar 0.32fF
C417 clk ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.32fF
C418 vdd cla_2/p0 0.43fF
C419 sumffo_2/ffo_0/nand_1/b cla_0/n 0.05fF
C420 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op nand_5/a 0.04fF
C421 ffo_0/nand_7/w_0_0# couto 0.04fF
C422 cinin ffipgarr_0/ffi_0/inv_0/w_0_6# 0.06fF
C423 y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.04fF
C424 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.06fF
C425 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C426 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C427 vdd nor_1/w_0_0# 0.15fF
C428 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_1/b 0.06fF
C429 clk sumffo_3/ffo_0/nand_3/b 0.33fF
C430 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.04fF
C431 vdd z1o 0.28fF
C432 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.04fF
C433 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C434 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_7/a 0.04fF
C435 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/nand_3/b 0.06fF
C436 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C437 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.45fF
C438 cla_1/inv_0/in gnd 0.35fF
C439 nor_4/b inv_9/in 0.16fF
C440 cla_0/n sumffo_2/ffo_0/nand_1/w_0_0# 0.13fF
C441 ffo_0/d ffo_0/inv_0/op 0.04fF
C442 sumffo_3/xor_0/inv_1/op sumffo_3/ffo_0/d 0.52fF
C443 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_0/b 0.13fF
C444 sumffo_2/xor_0/inv_1/w_0_6# vdd 0.06fF
C445 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_0/b 0.40fF
C446 vdd ffipgarr_0/ffi_0/nand_3/w_0_0# 0.11fF
C447 vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.34fF
C448 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.06fF
C449 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.06fF
C450 ffipgarr_0/ffipg_0/ffi_0/nand_3/a clk 0.13fF
C451 vdd cla_1/inv_0/w_0_6# 0.06fF
C452 inv_2/op nand_2/b 0.10fF
C453 vdd ffo_0/nand_6/w_0_0# 0.10fF
C454 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/op 1.63fF
C455 gnd cla_2/nor_1/w_0_0# 0.01fF
C456 gnd cla_1/nor_1/a_13_6# 0.01fF
C457 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C458 gnd sumffo_2/ffo_0/nand_3/a 0.03fF
C459 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C460 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_1/ffi_0/qbar 0.06fF
C461 gnd ffipgarr_0/ffipg_0/ffi_1/qbar 0.34fF
C462 gnd ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.10fF
C463 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.31fF
C464 sumffo_1/xor_0/inv_1/w_0_6# vdd 0.06fF
C465 vdd ffipgarr_0/ffi_0/nand_3/b 0.39fF
C466 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C467 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_0/op 0.08fF
C468 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.39fF
C469 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.31fF
C470 vdd sumffo_3/ffo_0/nand_1/a 0.30fF
C471 vdd ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.10fF
C472 sumffo_3/ffo_0/inv_0/w_0_6# gnd 0.01fF
C473 sumffo_1/ffo_0/nand_7/w_0_0# z2o 0.04fF
C474 clk ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# 0.06fF
C475 gnd ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.03fF
C476 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.04fF
C477 inv_7/op inv_8/w_0_6# 0.06fF
C478 cla_1/n nor_2/b 0.37fF
C479 sumffo_3/sbar vdd 0.28fF
C480 sumffo_2/xor_0/inv_0/op sumffo_2/ffo_0/d 0.06fF
C481 vdd ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# 0.10fF
C482 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C483 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.06fF
C484 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.06fF
C485 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C486 vdd sumffo_1/xor_0/inv_1/op 0.15fF
C487 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/d 0.04fF
C488 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C489 vdd nand_2/b 0.82fF
C490 cla_2/g1 cla_2/p1 0.00fF
C491 gnd ffipgarr_0/ffipg_0/ffi_1/nand_0/a_13_n26# 0.01fF
C492 vdd ffo_0/nand_7/w_0_0# 0.12fF
C493 vdd ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# 0.10fF
C494 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/w_n3_4# 0.06fF
C495 gnd sumffo_0/ffo_0/nand_0/b 0.38fF
C496 gnd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.00fF
C497 nor_0/b nand_5/a 2.65fF
C498 ffipgarr_0/ffipg_2/ffi_1/inv_0/op clk 0.32fF
C499 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.06fF
C500 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# y2in 0.06fF
C501 ffipgarr_0/ffipg_1/ffi_0/nand_6/a ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.04fF
C502 vdd ffo_0/nand_5/w_0_0# 0.10fF
C503 vdd sumffo_2/ffo_0/nand_6/a 0.30fF
C504 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.06fF
C505 gnd y2in 0.19fF
C506 inv_3/w_0_6# cla_1/l 0.06fF
C507 sumffo_2/ffo_0/nand_3/w_0_0# sumffo_2/ffo_0/nand_3/a 0.06fF
C508 gnd ffipgarr_0/ffi_0/nand_0/a_13_n26# 0.01fF
C509 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.33fF
C510 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.32fF
C511 ffipgarr_0/ffipg_1/ffi_0/inv_0/op clk 0.32fF
C512 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.04fF
C513 cla_1/g0 cla_0/inv_0/op 0.35fF
C514 sumffo_2/ffo_0/inv_1/w_0_6# sumffo_2/ffo_0/nand_0/b 0.03fF
C515 vdd z3o 0.28fF
C516 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C517 ffipgarr_0/ffipg_1/ffi_1/inv_1/op x2in 0.01fF
C518 sumffo_1/ffo_0/nand_5/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C519 gnd ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.03fF
C520 gnd cla_0/n 0.52fF
C521 cla_1/g0 cla_1/p0 1.76fF
C522 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.04fF
C523 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C524 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C525 nand_2/b cla_1/nor_0/w_0_0# 0.01fF
C526 sumffo_1/k cla_0/g0 0.07fF
C527 ffo_0/nand_7/a ffo_0/nand_1/b 0.13fF
C528 ffo_0/nand_1/w_0_0# ffo_0/nand_1/b 0.06fF
C529 vdd ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.10fF
C530 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.00fF
C531 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.13fF
C532 ffipgarr_0/ffipg_0/ffi_0/nand_1/b vdd 0.31fF
C533 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.32fF
C534 vdd inv_8/in 0.30fF
C535 cla_0/g0 cla_0/inv_0/in 0.16fF
C536 cla_2/inv_0/in cla_2/g0 0.16fF
C537 nor_4/a nor_4/b 0.35fF
C538 clk sumffo_1/ffo_0/nand_1/b 0.45fF
C539 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_3/a 0.06fF
C540 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# 0.06fF
C541 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/q 0.06fF
C542 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C543 vdd inv_4/op 0.25fF
C544 vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.34fF
C545 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.30fF
C546 vdd ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.10fF
C547 vdd ffipgarr_0/ffipg_3/ffi_1/qbar 0.33fF
C548 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C549 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C550 inv_6/in nor_3/w_0_0# 0.11fF
C551 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# gnd 0.00fF
C552 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.20fF
C553 cla_0/l cla_1/nand_0/w_0_0# 0.08fF
C554 vdd sumffo_3/k 0.31fF
C555 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C556 vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.10fF
C557 sumffo_3/xor_0/a_10_10# vdd 0.93fF
C558 vdd sumffo_3/ffo_0/nand_3/w_0_0# 0.11fF
C559 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_0/w_0_0# 0.04fF
C560 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C561 inv_3/w_0_6# gnd 0.01fF
C562 ffo_0/nand_3/a ffo_0/nand_3/w_0_0# 0.06fF
C563 ffo_0/nand_1/a ffo_0/nand_1/b 0.31fF
C564 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_1/b 0.13fF
C565 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/ffo_0/nand_7/a 0.06fF
C566 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/qbar 0.06fF
C567 cla_0/nor_0/a_13_6# nand_5/a 0.01fF
C568 vdd sumffo_3/xor_0/inv_1/w_0_6# 0.06fF
C569 sumffo_3/ffo_0/d sumffo_3/ffo_0/inv_0/op 0.04fF
C570 nand_5/a sumffo_0/xor_0/inv_0/op 0.20fF
C571 vdd cla_2/nand_0/w_0_0# 0.10fF
C572 clk ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.07fF
C573 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.30fF
C574 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_1/b 0.13fF
C575 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.06fF
C576 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# clk 0.06fF
C577 vdd ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.10fF
C578 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.06fF
C579 cla_1/p0 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C580 vdd ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.10fF
C581 vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.10fF
C582 sumffo_0/k vdd 0.31fF
C583 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.06fF
C584 gnd sumffo_2/ffo_0/nand_0/a_13_n26# 0.00fF
C585 gnd x3in 0.19fF
C586 clk sumffo_3/ffo_0/d 0.26fF
C587 sumffo_1/sbar z2o 0.32fF
C588 sumffo_1/ffo_0/nand_3/b clk 0.33fF
C589 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/sbar 0.04fF
C590 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/a 0.06fF
C591 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.06fF
C592 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.30fF
C593 gnd y3in 0.19fF
C594 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.13fF
C595 vdd ffipgarr_0/ffipg_1/ffi_1/q 1.33fF
C596 vdd ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.10fF
C597 cla_1/inv_0/op cla_1/inv_0/in 0.04fF
C598 inv_1/w_0_6# nand_5/a 0.06fF
C599 ffo_0/nand_3/b ffo_0/nand_1/b 0.32fF
C600 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_3/a 0.13fF
C601 nor_0/a nor_0/w_0_0# 0.06fF
C602 ffo_0/d vdd 0.19fF
C603 x4in ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.01fF
C604 vdd ffipgarr_0/ffi_0/nand_1/b 0.31fF
C605 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# 0.06fF
C606 sumffo_0/ffo_0/nand_4/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C607 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.06fF
C608 gnd ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.26fF
C609 cla_1/g0 gnd 0.76fF
C610 gnd inv_6/in 0.24fF
C611 gnd sumffo_3/ffo_0/nand_1/b 0.26fF
C612 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.04fF
C613 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.04fF
C614 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.13fF
C615 vdd sumffo_1/ffo_0/inv_0/op 0.17fF
C616 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/inv_0/w_0_6# 0.03fF
C617 sumffo_0/ffo_0/nand_6/w_0_0# vdd 0.10fF
C618 vdd ffipgarr_0/ffipg_2/ffi_0/q 0.38fF
C619 ffipgarr_0/ffipg_0/ffi_0/nand_3/a ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.04fF
C620 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C621 vdd sumffo_0/ffo_0/nand_2/w_0_0# 0.10fF
C622 ffo_0/nand_0/w_0_0# ffo_0/nand_1/a 0.04fF
C623 ffipgarr_0/ffipg_0/ffi_1/inv_0/op gnd 0.10fF
C624 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C625 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_7/a 0.13fF
C626 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.39fF
C627 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C628 gnd inv_0/in 0.24fF
C629 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C630 cla_2/l cla_0/n 0.31fF
C631 sumffo_3/ffo_0/d sumffo_3/ffo_0/nand_0/b 0.40fF
C632 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/b 0.06fF
C633 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.33fF
C634 ffipgarr_0/ffi_0/inv_1/op ffipgarr_0/ffi_0/nand_6/a 0.13fF
C635 gnd ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.22fF
C636 gnd inv_3/in 0.36fF
C637 vdd ffipgarr_0/ffipg_0/ffi_1/q 1.35fF
C638 clk ffipgarr_0/ffi_0/nand_0/w_0_0# 0.06fF
C639 vdd nor_2/b 0.35fF
C640 sumffo_1/sbar sumffo_1/ffo_0/nand_6/a 0.00fF
C641 gnd cla_2/p1 0.69fF
C642 sumffo_2/k cla_1/g0 0.56fF
C643 gnd sumffo_2/sbar 0.34fF
C644 cla_2/p1 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C645 cla_1/p0 ffipgarr_0/ffipg_1/ffi_0/q 0.21fF
C646 sumffo_0/xor_0/w_n3_4# vdd 0.12fF
C647 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_3/b 0.00fF
C648 ffipgarr_0/ffi_0/nand_3/a ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C649 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.30fF
C650 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.30fF
C651 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.06fF
C652 inv_5/in inv_5/w_0_6# 0.10fF
C653 z1o sumffo_0/ffo_0/nand_6/a 0.31fF
C654 gnd z2o 0.52fF
C655 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.20fF
C656 sumffo_0/ffo_0/nand_7/w_0_0# sumffo_0/sbar 0.06fF
C657 ffipgarr_0/ffipg_3/ffi_0/nand_6/a ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.06fF
C658 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.31fF
C659 gnd inv_1/in 0.22fF
C660 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/sbar 0.06fF
C661 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C662 sumffo_3/xor_0/inv_1/op inv_4/op 0.22fF
C663 sumffo_3/ffo_0/nand_7/w_0_0# sumffo_3/ffo_0/nand_7/a 0.06fF
C664 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C665 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/a 0.31fF
C666 cla_0/nor_1/w_0_0# cla_0/inv_0/in 0.05fF
C667 cla_0/l cla_1/n 0.18fF
C668 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op sumffo_3/k 0.06fF
C669 gnd ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.26fF
C670 inv_8/in nor_4/b 0.04fF
C671 inv_4/op inv_4/in 0.04fF
C672 clk ffo_0/nand_0/b 0.04fF
C673 sumffo_3/xor_0/inv_1/op sumffo_3/k 0.06fF
C674 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/w_0_0# 0.04fF
C675 vdd sumffo_0/ffo_0/nand_7/w_0_0# 0.10fF
C676 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.00fF
C677 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.31fF
C678 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# y2in 0.06fF
C679 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/qbar 0.00fF
C680 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/ffi_1/q 0.27fF
C681 ffipgarr_0/ffipg_0/ffi_0/q nand_2/b 0.90fF
C682 vdd inv_5/w_0_6# 0.15fF
C683 gnd x1in 0.19fF
C684 sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/inv_1/w_0_6# 0.03fF
C685 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.31fF
C686 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/qbar 0.32fF
C687 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.06fF
C688 vdd cla_1/nand_0/w_0_0# 0.10fF
C689 cla_0/inv_0/op cla_0/inv_0/in 0.04fF
C690 cla_1/g0 ffipgarr_0/ffipg_2/ffi_1/q 0.93fF
C691 nor_1/b cla_0/l 0.10fF
C692 inv_7/op inv_7/w_0_6# 0.03fF
C693 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_7/w_0_0# 0.06fF
C694 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.52fF
C695 nor_0/a inv_0/in 0.02fF
C696 gnd sumffo_1/ffo_0/nand_6/a 0.03fF
C697 gnd sumffo_2/ffo_0/nand_7/a 0.03fF
C698 cla_2/g1 ffipgarr_0/ffipg_3/ffi_0/q 0.13fF
C699 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.04fF
C700 vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.10fF
C701 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/q 0.00fF
C702 sumffo_1/k cla_1/p0 0.05fF
C703 sumffo_1/xor_0/w_n3_4# sumffo_1/ffo_0/d 0.02fF
C704 vdd cla_2/n 0.28fF
C705 vdd ffipgarr_0/ffi_0/inv_0/op 0.17fF
C706 vdd ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.10fF
C707 ffipgarr_0/ffipg_1/ffi_1/inv_1/op clk 0.07fF
C708 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.13fF
C709 cla_1/p0 cla_0/inv_0/in 0.02fF
C710 cla_0/nor_1/a_13_6# gnd 0.01fF
C711 cla_2/g1 cla_2/g0 0.13fF
C712 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C713 gnd ffipgarr_0/ffipg_3/ffi_0/qbar 0.34fF
C714 gnd ffipgarr_0/ffipg_1/ffi_0/q 2.58fF
C715 nand_5/a inv_8/in 0.00fF
C716 sumffo_0/xor_0/a_10_10# vdd 0.93fF
C717 vdd ffipgarr_0/ffi_0/nand_7/w_0_0# 0.10fF
C718 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.06fF
C719 cla_0/n sumffo_2/ffo_0/nand_3/a 0.07fF
C720 gnd ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.03fF
C721 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op sumffo_3/k 0.52fF
C722 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C723 sumffo_2/ffo_0/nand_7/w_0_0# sumffo_2/ffo_0/nand_7/a 0.06fF
C724 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# 0.04fF
C725 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C726 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.45fF
C727 vdd sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C728 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_7/a 0.13fF
C729 cla_2/l cla_2/p1 0.02fF
C730 gnd y4in 0.19fF
C731 gnd ffipgarr_0/ffi_0/nand_6/a 0.03fF
C732 gnd ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.34fF
C733 ffo_0/nand_5/w_0_0# clk 0.06fF
C734 sumffo_3/sbar z4o 0.32fF
C735 clk sumffo_2/ffo_0/nand_6/a 0.13fF
C736 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.00fF
C737 vdd ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.10fF
C738 ffipgarr_0/ffipg_2/ffi_0/inv_0/op ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.03fF
C739 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.06fF
C740 vdd cla_0/nor_0/w_0_0# 0.32fF
C741 vdd inv_7/in 0.34fF
C742 vdd sumffo_3/ffo_0/nand_7/a 0.30fF
C743 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.06fF
C744 gnd sumffo_3/ffo_0/nand_6/a 0.03fF
C745 gnd ffipgarr_0/ffipg_1/ffi_1/nand_0/a_13_n26# 0.01fF
C746 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.13fF
C747 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/b 0.13fF
C748 vdd sumffo_1/ffo_0/nand_1/a 0.30fF
C749 sumffo_0/k nand_5/a 0.41fF
C750 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.75fF
C751 ffipgarr_0/ffi_0/nand_7/a ffipgarr_0/ffi_0/nand_5/w_0_0# 0.04fF
C752 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C753 vdd cla_2/inv_0/w_0_6# 0.06fF
C754 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# 0.10fF
C755 sumffo_0/k ffipgarr_0/ffipg_0/ffi_0/q 0.07fF
C756 vdd ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# 0.10fF
C757 nor_2/b inv_4/in 0.16fF
C758 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/b 0.31fF
C759 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# 0.06fF
C760 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C761 vdd cla_2/nor_0/w_0_0# 0.31fF
C762 gnd x4in 0.19fF
C763 clk ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C764 vdd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.10fF
C765 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.13fF
C766 sumffo_1/k gnd 0.35fF
C767 cla_1/g0 cla_1/inv_0/in 0.16fF
C768 cla_0/inv_0/in gnd 0.35fF
C769 vdd sumffo_2/ffo_0/nand_4/w_0_0# 0.10fF
C770 vdd ffipgarr_0/ffi_0/nand_5/w_0_0# 0.10fF
C771 vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.10fF
C772 gnd ffo_0/nand_1/b 0.26fF
C773 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.04fF
C774 inv_0/op cla_0/g0 0.32fF
C775 vdd ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# 0.10fF
C776 gnd sumffo_3/ffo_0/nand_3/a 0.03fF
C777 sumffo_1/ffo_0/nand_0/w_0_0# sumffo_1/ffo_0/nand_0/b 0.06fF
C778 sumffo_0/ffo_0/inv_1/w_0_6# sumffo_0/ffo_0/nand_0/b 0.03fF
C779 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C780 ffipgarr_0/ffipg_0/ffi_1/inv_0/op ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.03fF
C781 ffipgarr_0/ffipg_0/ffi_1/nand_1/a clk 0.13fF
C782 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.06fF
C783 inv_2/op cla_0/l 0.06fF
C784 vdd sumffo_1/ffo_0/nand_4/w_0_0# 0.10fF
C785 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.30fF
C786 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.30fF
C787 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C788 sumffo_3/ffo_0/nand_6/a sumffo_3/ffo_0/nand_4/w_0_0# 0.04fF
C789 gnd ffipgarr_0/ffipg_3/ffi_1/inv_0/op 0.10fF
C790 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C791 vdd cla_1/n 0.28fF
C792 vdd cla_0/inv_0/w_0_6# 0.06fF
C793 ffo_0/nand_6/a couto 0.31fF
C794 sumffo_0/ffo_0/nand_6/w_0_0# sumffo_0/ffo_0/nand_6/a 0.06fF
C795 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.30fF
C796 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/w_0_0# 0.04fF
C797 inv_3/w_0_6# cla_0/n 0.00fF
C798 ffipgarr_0/ffipg_0/ffi_1/q nand_5/a 0.02fF
C799 inv_2/in nor_1/w_0_0# 0.11fF
C800 gnd sumffo_3/ffo_0/nand_3/b 0.35fF
C801 clk ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.13fF
C802 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/qbar 0.31fF
C803 vdd ffo_0/inv_0/op 0.17fF
C804 vdd sumffo_1/xor_0/w_n3_4# 0.12fF
C805 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.32fF
C806 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_1/q 0.73fF
C807 vdd cla_0/l 1.74fF
C808 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.04fF
C809 gnd sumffo_1/ffo_0/nand_0/w_0_0# 0.08fF
C810 gnd ffipgarr_0/ffipg_1/ffi_0/qbar 0.34fF
C811 cla_2/p1 cla_2/nor_1/w_0_0# 0.06fF
C812 nor_1/b vdd 0.35fF
C813 ffo_0/nand_0/b ffo_0/nand_1/a 0.13fF
C814 sumffo_0/xor_0/w_n3_4# nand_5/a 0.06fF
C815 sumffo_0/ffo_0/nand_7/a sumffo_0/sbar 0.31fF
C816 ffipgarr_0/ffipg_3/ffi_1/nand_3/a ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.04fF
C817 gnd ffipgarr_0/ffipg_3/ffi_1/q 0.93fF
C818 clk ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.13fF
C819 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# clk 0.06fF
C820 ffipgarr_0/ffipg_0/ffi_0/nand_3/a gnd 0.03fF
C821 vdd sumffo_3/ffo_0/nand_6/w_0_0# 0.10fF
C822 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C823 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.31fF
C824 vdd sumffo_1/ffo_0/d 0.04fF
C825 vdd sumffo_0/ffo_0/nand_1/b 0.31fF
C826 gnd ffipgarr_0/ffipg_3/ffi_0/q 2.62fF
C827 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/q 0.31fF
C828 cla_1/g0 cla_0/n 0.13fF
C829 vdd sumffo_0/ffo_0/nand_7/a 0.30fF
C830 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.31fF
C831 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.31fF
C832 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.33fF
C833 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# 0.06fF
C834 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C835 sumffo_1/k nor_0/a 0.06fF
C836 vdd sumffo_0/ffo_0/nand_0/w_0_0# 0.10fF
C837 gnd ffipgarr_0/ffipg_2/ffi_1/qbar 0.34fF
C838 gnd cla_2/g0 0.32fF
C839 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C840 x1in ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C841 inv_7/op inv_8/in 0.13fF
C842 inv_0/in nor_0/w_0_0# 0.11fF
C843 ffo_0/nand_7/a ffo_0/nand_7/w_0_0# 0.06fF
C844 vdd ffo_0/nand_6/a 0.30fF
C845 vdd sumffo_3/ffo_0/nand_7/w_0_0# 0.10fF
C846 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C847 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_2/w_0_0# 0.06fF
C848 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# ffipgarr_0/ffipg_0/ffi_1/qbar 0.06fF
C849 cla_0/g0 nand_2/b 1.01fF
C850 ffo_0/nand_7/a ffo_0/nand_5/w_0_0# 0.04fF
C851 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C852 vdd ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.10fF
C853 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.31fF
C854 gnd ffipgarr_0/ffipg_2/ffi_1/inv_0/op 0.10fF
C855 gnd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C856 vdd ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# 0.10fF
C857 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.06fF
C858 ffipgarr_0/ffipg_1/ffi_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.03fF
C859 vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C860 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.04fF
C861 inv_3/in cla_0/n 0.02fF
C862 vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.34fF
C863 vdd ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.34fF
C864 gnd ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.10fF
C865 sumffo_2/xor_0/inv_0/op gnd 0.17fF
C866 ffipgarr_0/ffipg_1/ffi_0/nand_1/a clk 0.13fF
C867 vdd ffipgarr_0/ffipg_0/ffi_1/inv_1/op 1.63fF
C868 ffipgarr_0/ffipg_0/ffi_1/nand_3/a clk 0.13fF
C869 ffipgarr_0/ffipg_0/ffi_1/nand_1/b gnd 0.26fF
C870 ffipgarr_0/ffipg_0/ffi_0/nand_1/a ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.00fF
C871 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C872 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.30fF
C873 nand_2/b cla_0/nand_0/w_0_0# 0.01fF
C874 vdd couto 0.28fF
C875 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.06fF
C876 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.04fF
C877 sumffo_0/xor_0/a_10_10# nand_5/a 0.12fF
C878 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.03fF
C879 nand_5/a ffipgarr_0/ffi_0/nand_7/w_0_0# 0.04fF
C880 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.15fF
C881 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.06fF
C882 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# 0.11fF
C883 cla_2/inv_0/op cla_2/inv_0/w_0_6# 0.03fF
C884 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.33fF
C885 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_2/w_0_0# 0.06fF
C886 ffipgarr_0/ffipg_3/ffi_1/inv_1/op ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C887 vdd ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.10fF
C888 gnd sumffo_1/ffo_0/nand_1/b 0.26fF
C889 gnd ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.35fF
C890 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.06fF
C891 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_1/w_0_0# 0.04fF
C892 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# 0.06fF
C893 gnd ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.35fF
C894 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# 0.04fF
C895 inv_3/w_0_6# inv_3/in 0.10fF
C896 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.06fF
C897 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/inv_0/op 0.06fF
C898 vdd inv_5/in 0.30fF
C899 vdd sumffo_1/ffo_0/nand_6/w_0_0# 0.10fF
C900 vdd inv_2/op 0.34fF
C901 vdd sumffo_0/ffo_0/nand_3/w_0_0# 0.11fF
C902 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C903 cla_0/nor_0/w_0_0# nand_5/a 0.01fF
C904 gnd inv_9/in 0.24fF
C905 gnd nor_0/b 0.59fF
C906 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.04fF
C907 cla_1/n inv_4/in 0.02fF
C908 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/w_0_0# 0.04fF
C909 inv_2/op sumffo_2/xor_0/inv_1/op 0.22fF
C910 sumffo_2/k sumffo_2/xor_0/inv_0/op 0.27fF
C911 sumffo_2/ffo_0/nand_3/a sumffo_2/ffo_0/nand_2/w_0_0# 0.04fF
C912 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_0/op 0.08fF
C913 vdd sumffo_0/sbar 0.28fF
C914 vdd ffipgarr_0/ffi_0/nand_7/a 0.30fF
C915 vdd ffipgarr_0/ffi_0/nand_4/w_0_0# 0.10fF
C916 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.75fF
C917 vdd ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# 0.11fF
C918 ffipgarr_0/ffipg_2/ffi_0/inv_1/op y3in 0.01fF
C919 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C920 gnd ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.22fF
C921 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C922 vdd ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# 0.10fF
C923 ffo_0/nand_2/w_0_0# ffo_0/nand_3/a 0.04fF
C924 ffipgarr_0/ffi_0/inv_0/op clk 0.32fF
C925 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_3/b 0.00fF
C926 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.30fF
C927 vdd ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.39fF
C928 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_0/q 0.06fF
C929 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/qbar 0.32fF
C930 cla_0/g0 ffipgarr_0/ffipg_1/ffi_1/q 0.84fF
C931 gnd sumffo_3/ffo_0/d 0.37fF
C932 sumffo_1/ffo_0/nand_3/b gnd 0.35fF
C933 ffipgarr_0/ffi_0/nand_6/w_0_0# ffipgarr_0/ffi_0/nand_6/a 0.06fF
C934 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# 0.06fF
C935 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# clk 0.06fF
C936 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_3/b 0.00fF
C937 nor_3/b inv_5/w_0_6# 0.03fF
C938 nor_3/w_0_0# nor_4/a 0.03fF
C939 vdd sumffo_2/xor_0/inv_1/op 0.15fF
C940 sumffo_0/ffo_0/d sumffo_0/xor_0/inv_0/op 0.06fF
C941 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.11fF
C942 ffipgarr_0/ffipg_2/ffi_0/nand_7/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.31fF
C943 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.04fF
C944 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.06fF
C945 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C946 gnd cla_1/nor_1/w_0_0# 0.01fF
C947 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C948 cla_1/p0 cla_2/p0 0.24fF
C949 clk sumffo_1/ffo_0/inv_1/w_0_6# 0.06fF
C950 vdd ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.10fF
C951 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/inv_1/op 0.33fF
C952 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/nand_0/w_0_0# 0.06fF
C953 gnd sumffo_0/ffo_0/nand_1/a 0.03fF
C954 cla_1/inv_0/op cla_2/g0 0.35fF
C955 cla_0/n sumffo_2/ffo_0/nand_2/w_0_0# 0.13fF
C956 nor_3/b cla_2/n 0.37fF
C957 ffo_0/nand_3/a ffo_0/nand_0/b 0.13fF
C958 sumffo_0/ffo_0/nand_3/b sumffo_0/ffo_0/nand_3/a 0.31fF
C959 vdd ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# 0.10fF
C960 gnd ffipgarr_0/ffipg_1/ffi_0/nand_3/b 0.35fF
C961 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.20fF
C962 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C963 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_1/nand_1/a 0.04fF
C964 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_0/ffi_0/inv_1/op 0.06fF
C965 cla_2/p0 cla_1/l 0.02fF
C966 cla_0/l sumffo_2/ffo_0/nand_0/w_0_0# 0.17fF
C967 cla_0/nor_1/w_0_0# nand_2/b 0.02fF
C968 inv_4/op nor_2/w_0_0# 0.03fF
C969 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C970 vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C971 vdd ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.15fF
C972 vdd cla_1/nor_0/w_0_0# 0.32fF
C973 inv_2/op sumffo_2/xor_0/a_10_10# 0.12fF
C974 gnd ffo_0/nand_2/w_0_0# 0.00fF
C975 gnd sumffo_0/xor_0/inv_0/op 0.17fF
C976 gnd ffipgarr_0/ffi_0/nand_0/w_0_0# 0.00fF
C977 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.04fF
C978 cla_0/l nand_5/a 0.36fF
C979 nor_0/a nor_0/b 0.39fF
C980 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/q 0.06fF
C981 vdd x2in 0.04fF
C982 sumffo_3/ffo_0/nand_7/a z4o 0.00fF
C983 gnd nor_4/a 0.15fF
C984 inv_1/w_0_6# gnd 0.01fF
C985 gnd sumffo_0/ffo_0/nand_3/a 0.03fF
C986 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.04fF
C987 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# clk 0.06fF
C988 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C989 clk sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C990 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C991 vdd ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.34fF
C992 ffipgarr_0/ffipg_0/ffi_1/inv_0/op x1in 0.04fF
C993 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# 0.12fF
C994 vdd sumffo_2/xor_0/a_10_10# 0.93fF
C995 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C996 inv_0/op gnd 0.10fF
C997 cla_0/l cla_1/nand_0/a_13_n26# 0.01fF
C998 cla_1/g0 ffipgarr_0/ffipg_1/ffi_0/q 0.29fF
C999 cla_1/inv_0/in cla_2/g0 0.04fF
C1000 sumffo_1/ffo_0/nand_3/a sumffo_1/ffo_0/nand_2/w_0_0# 0.04fF
C1001 gnd ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.03fF
C1002 nand_2/b cla_1/p0 2.00fF
C1003 clk sumffo_1/ffo_0/nand_4/w_0_0# 0.06fF
C1004 clk ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.13fF
C1005 ffipgarr_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffi_0/nand_1/b 0.06fF
C1006 vdd ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# 0.10fF
C1007 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.00fF
C1008 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# ffipgarr_0/ffipg_2/ffi_0/qbar 0.06fF
C1009 ffipgarr_0/ffipg_1/ffi_1/nand_1/a clk 0.13fF
C1010 sumffo_0/ffo_0/nand_7/a sumffo_0/ffo_0/nand_5/w_0_0# 0.04fF
C1011 ffipgarr_0/ffipg_3/ffi_1/nand_1/a ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.00fF
C1012 vdd ffipgarr_0/ffipg_2/ffi_0/qbar 0.33fF
C1013 cla_2/g0 cla_2/nor_1/w_0_0# 0.06fF
C1014 gnd ffo_0/nand_0/b 0.43fF
C1015 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/a 0.31fF
C1016 cla_2/nand_0/w_0_0# cla_2/g1 0.06fF
C1017 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.06fF
C1018 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# 0.06fF
C1019 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.45fF
C1020 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C1021 cla_2/p0 gnd 0.74fF
C1022 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/nand_3/a 0.04fF
C1023 vdd sumffo_1/xor_0/inv_0/w_0_6# 0.09fF
C1024 clk ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.13fF
C1025 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.04fF
C1026 x2in ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.06fF
C1027 nand_2/b cla_1/l 0.35fF
C1028 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_1/b 0.06fF
C1029 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.04fF
C1030 cla_0/l clk 0.12fF
C1031 z1o gnd 0.52fF
C1032 cla_2/inv_0/in cla_2/inv_0/w_0_6# 0.06fF
C1033 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.15fF
C1034 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.04fF
C1035 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.00fF
C1036 vdd ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.34fF
C1037 vdd sumffo_3/xor_0/inv_1/op 0.15fF
C1038 sumffo_2/sbar sumffo_2/ffo_0/nand_7/a 0.31fF
C1039 vdd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.06fF
C1040 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.06fF
C1041 inv_7/op inv_7/in 0.04fF
C1042 gnd ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.03fF
C1043 z2o sumffo_1/ffo_0/nand_6/a 0.31fF
C1044 vdd ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.34fF
C1045 ffipgarr_0/ffipg_2/ffi_1/inv_1/op ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.04fF
C1046 gnd ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.22fF
C1047 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/q 0.06fF
C1048 vdd sumffo_0/ffo_0/inv_0/op 0.17fF
C1049 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/ffi_0/q 0.12fF
C1050 clk sumffo_1/ffo_0/d 0.05fF
C1051 vdd inv_4/in 0.09fF
C1052 clk sumffo_0/ffo_0/nand_1/b 0.45fF
C1053 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.31fF
C1054 nor_2/b nor_2/w_0_0# 0.06fF
C1055 cla_2/l inv_7/w_0_6# 0.06fF
C1056 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.35fF
C1057 gnd ffipgarr_0/ffi_0/nand_3/b 0.35fF
C1058 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/qbar 0.32fF
C1059 sumffo_3/ffo_0/nand_1/a gnd 0.03fF
C1060 sumffo_1/ffo_0/nand_3/w_0_0# sumffo_1/ffo_0/nand_1/b 0.04fF
C1061 vdd cla_2/inv_0/op 0.17fF
C1062 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.00fF
C1063 sumffo_2/k cla_2/p0 0.05fF
C1064 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.75fF
C1065 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# clk 0.06fF
C1066 vdd nor_4/b 0.41fF
C1067 sumffo_1/ffo_0/nand_1/w_0_0# sumffo_1/ffo_0/nand_1/a 0.06fF
C1068 sumffo_3/ffo_0/nand_6/w_0_0# z4o 0.06fF
C1069 ffipgarr_0/ffi_0/nand_1/b ffipgarr_0/ffi_0/inv_1/op 0.45fF
C1070 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C1071 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C1072 cla_1/g0 cla_0/inv_0/in 0.04fF
C1073 sumffo_3/sbar gnd 0.34fF
C1074 clk ffo_0/nand_6/a 0.13fF
C1075 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C1076 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C1077 gnd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.17fF
C1078 nand_2/b gnd 1.54fF
C1079 vdd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.15fF
C1080 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# nand_5/a 0.02fF
C1081 clk ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# 0.06fF
C1082 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C1083 gnd sumffo_2/ffo_0/nand_6/a 0.03fF
C1084 ffipgarr_0/ffi_0/nand_7/a nand_5/a 0.00fF
C1085 ffipgarr_0/ffipg_1/ffi_0/inv_0/op y2in 0.04fF
C1086 cla_0/l sumffo_2/ffo_0/nand_1/a 0.15fF
C1087 sumffo_3/ffo_0/nand_7/w_0_0# z4o 0.04fF
C1088 sumffo_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C1089 vdd sumffo_2/ffo_0/nand_0/w_0_0# 0.10fF
C1090 vdd ffipgarr_0/ffi_0/nand_1/a 0.30fF
C1091 ffo_0/nand_3/w_0_0# ffo_0/nand_1/b 0.04fF
C1092 gnd z3o 0.52fF
C1093 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.06fF
C1094 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.00fF
C1095 ffipgarr_0/ffipg_1/ffi_1/q cla_1/p0 0.22fF
C1096 ffipgarr_0/ffipg_0/ffi_1/inv_1/op clk 0.07fF
C1097 ffipgarr_0/ffipg_0/ffi_0/nand_1/a clk 0.13fF
C1098 ffo_0/qbar ffo_0/nand_6/w_0_0# 0.04fF
C1099 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_3/w_0_0# 0.06fF
C1100 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# cla_0/g0 0.04fF
C1101 vdd nand_5/a 1.48fF
C1102 sumffo_0/sbar sumffo_0/ffo_0/nand_6/a 0.00fF
C1103 ffo_0/d ffo_0/inv_0/w_0_6# 0.06fF
C1104 vdd sumffo_0/ffo_0/nand_5/w_0_0# 0.10fF
C1105 vdd ffipgarr_0/ffi_0/nand_3/a 0.30fF
C1106 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C1107 vdd ffipgarr_0/ffipg_0/ffi_0/q 0.38fF
C1108 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_1/b 0.32fF
C1109 cla_2/l cla_2/p0 0.16fF
C1110 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.32fF
C1111 cla_2/p0 ffipgarr_0/ffipg_2/ffi_1/q 0.22fF
C1112 ffipgarr_0/ffipg_0/ffi_0/nand_1/b gnd 0.26fF
C1113 gnd inv_8/in 0.13fF
C1114 sumffo_2/k nand_2/b 0.03fF
C1115 sumffo_2/ffo_0/nand_7/w_0_0# z3o 0.04fF
C1116 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.31fF
C1117 clk ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# 0.06fF
C1118 ffipgarr_0/ffi_0/nand_6/w_0_0# nor_0/b 0.04fF
C1119 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.06fF
C1120 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/nor_0/a_13_6# 0.01fF
C1121 ffipgarr_0/ffipg_1/ffi_0/nand_3/a ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.06fF
C1122 vdd ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# 0.11fF
C1123 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C1124 vdd sumffo_0/ffo_0/nand_6/a 0.30fF
C1125 vdd ffipgarr_0/ffipg_0/ffi_0/inv_1/op 1.63fF
C1126 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.33fF
C1127 gnd inv_4/op 0.21fF
C1128 ffipgarr_0/ffipg_3/ffi_1/nand_1/b ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.32fF
C1129 gnd ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.03fF
C1130 ffipgarr_0/ffipg_0/ffi_1/nand_1/a gnd 0.15fF
C1131 sumffo_3/ffo_0/inv_0/w_0_6# sumffo_3/ffo_0/d 0.06fF
C1132 vdd sumffo_2/ffo_0/d 0.04fF
C1133 vdd ffipgarr_0/ffipg_2/ffi_1/inv_1/op 1.63fF
C1134 gnd ffipgarr_0/ffipg_3/ffi_1/qbar 0.34fF
C1135 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# y3in 0.06fF
C1136 inv_2/op clk 1.02fF
C1137 nor_0/b nor_0/w_0_0# 0.06fF
C1138 vdd sumffo_0/ffo_0/nand_1/w_0_0# 0.10fF
C1139 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.93fF
C1140 ffo_0/qbar ffo_0/nand_7/w_0_0# 0.06fF
C1141 sumffo_2/xor_0/inv_1/op sumffo_2/ffo_0/d 0.52fF
C1142 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.06fF
C1143 gnd sumffo_3/k 0.35fF
C1144 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/a 0.00fF
C1145 cla_1/g0 cla_2/g0 0.13fF
C1146 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op nand_5/a 0.04fF
C1147 vdd sumffo_1/ffo_0/nand_5/w_0_0# 0.10fF
C1148 sumffo_0/ffo_0/d sumffo_0/ffo_0/nand_2/w_0_0# 0.06fF
C1149 cla_2/g1 cla_2/n 0.13fF
C1150 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C1151 ffipgarr_0/ffipg_2/ffi_1/inv_0/op x3in 0.04fF
C1152 nand_2/b nor_0/a 1.53fF
C1153 vdd sumffo_3/ffo_0/inv_0/op 0.17fF
C1154 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/b 0.32fF
C1155 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op 0.20fF
C1156 cla_2/nand_0/w_0_0# gnd 0.01fF
C1157 gnd ffipgarr_0/ffipg_3/ffi_0/nand_3/a 0.03fF
C1158 sumffo_0/xor_0/w_n3_4# sumffo_0/xor_0/inv_1/op 0.06fF
C1159 vdd ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# 0.10fF
C1160 vdd ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.34fF
C1161 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C1162 vdd ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1163 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# 0.04fF
C1164 sumffo_0/k gnd 0.41fF
C1165 cla_2/p1 ffipgarr_0/ffipg_3/ffi_1/q 0.22fF
C1166 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_4/w_0_0# 0.06fF
C1167 ffipgarr_0/ffipg_1/ffi_0/nand_3/a clk 0.13fF
C1168 vdd clk 12.15fF
C1169 nor_1/b inv_2/in 0.16fF
C1170 gnd ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.03fF
C1171 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_1/qbar 0.04fF
C1172 ffipgarr_0/ffipg_1/ffi_1/q gnd 0.93fF
C1173 nand_2/b ffipgarr_0/ffipg_2/ffi_1/q 0.69fF
C1174 nor_3/b inv_5/in 0.04fF
C1175 ffo_0/d gnd 0.26fF
C1176 y4in ffipgarr_0/ffipg_3/ffi_0/inv_0/op 0.04fF
C1177 cla_2/p1 ffipgarr_0/ffipg_3/ffi_0/q 0.03fF
C1178 gnd ffipgarr_0/ffi_0/nand_1/b 0.26fF
C1179 cla_1/inv_0/op cla_1/inv_0/w_0_6# 0.03fF
C1180 nor_4/w_0_0# inv_9/in 0.11fF
C1181 sumffo_1/k ffipgarr_0/ffipg_1/ffi_0/q 0.07fF
C1182 sumffo_3/ffo_0/nand_5/w_0_0# sumffo_3/ffo_0/nand_7/a 0.04fF
C1183 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/w_0_0# 0.06fF
C1184 sumffo_0/ffo_0/nand_1/a sumffo_0/ffo_0/nand_0/b 0.13fF
C1185 cla_2/p0 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C1186 vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.10fF
C1187 vdd z4o 0.28fF
C1188 cla_2/g0 cla_2/p1 0.30fF
C1189 sumffo_3/ffo_0/nand_2/w_0_0# sumffo_3/ffo_0/d 0.06fF
C1190 sumffo_1/ffo_0/inv_0/op gnd 0.10fF
C1191 sumffo_0/xor_0/w_n3_4# sumffo_0/ffo_0/d 0.02fF
C1192 gnd ffipgarr_0/ffipg_2/ffi_0/q 2.62fF
C1193 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.04fF
C1194 clk ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# 0.06fF
C1195 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C1196 cla_0/l cla_0/nand_0/w_0_0# 0.15fF
C1197 vdd sumffo_1/ffo_0/nand_7/a 0.30fF
C1198 vdd ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1199 cla_2/p0 cla_1/inv_0/in 0.02fF
C1200 ffipgarr_0/ffipg_1/ffi_1/inv_1/op ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.33fF
C1201 gnd ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.35fF
C1202 nor_3/b vdd 0.35fF
C1203 vdd sumffo_3/ffo_0/nand_0/b 0.15fF
C1204 sumffo_2/ffo_0/d sumffo_2/xor_0/a_10_10# 0.45fF
C1205 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C1206 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# 0.06fF
C1207 sumffo_0/ffo_0/nand_0/b sumffo_0/ffo_0/nand_3/a 0.13fF
C1208 gnd ffipgarr_0/ffipg_0/ffi_1/q 0.94fF
C1209 gnd nor_2/b 0.10fF
C1210 vdd cla_2/inv_0/in 0.05fF
C1211 x4in ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.06fF
C1212 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.39fF
C1213 x2in clk 0.70fF
C1214 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.31fF
C1215 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C1216 cla_1/n nor_2/w_0_0# 0.06fF
C1217 ffo_0/nand_7/a couto 0.00fF
C1218 vdd sumffo_2/ffo_0/nand_1/a 0.30fF
C1219 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/a 0.31fF
C1220 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/qbar 0.32fF
C1221 gnd ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.14fF
C1222 gnd ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.03fF
C1223 sumffo_2/k ffipgarr_0/ffipg_2/ffi_0/q 0.07fF
C1224 inv_0/op nor_0/w_0_0# 0.03fF
C1225 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.04fF
C1226 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.31fF
C1227 ffipgarr_0/ffipg_0/ffi_0/inv_1/op ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.13fF
C1228 sumffo_0/k nor_0/a 0.05fF
C1229 nor_3/w_0_0# cla_2/n 0.06fF
C1230 vdd inv_7/op 0.15fF
C1231 inv_0/in nor_0/b 0.16fF
C1232 ffipgarr_0/ffipg_3/ffi_1/inv_0/op ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# 0.03fF
C1233 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/qbar 0.32fF
C1234 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/qbar 0.00fF
C1235 vdd ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.17fF
C1236 vdd sumffo_1/ffo_0/nand_1/w_0_0# 0.10fF
C1237 vdd sumffo_2/xor_0/inv_0/w_0_6# 0.09fF
C1238 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.00fF
C1239 ffipgarr_0/ffi_0/nand_5/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C1240 y3in ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# 0.06fF
C1241 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.13fF
C1242 sumffo_0/xor_0/a_10_10# sumffo_0/ffo_0/d 0.45fF
C1243 ffipgarr_0/ffipg_3/ffi_0/nand_3/a ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.06fF
C1244 nor_4/a nor_4/w_0_0# 0.06fF
C1245 cla_0/nor_0/w_0_0# cla_1/p0 0.06fF
C1246 gnd inv_5/w_0_6# 0.01fF
C1247 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.06fF
C1248 ffipgarr_0/ffi_0/inv_0/op cinin 0.04fF
C1249 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# 0.06fF
C1250 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C1251 inv_2/op inv_2/in 0.04fF
C1252 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/a 0.04fF
C1253 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/inv_0/w_0_6# 0.03fF
C1254 ffipgarr_0/ffipg_3/ffi_1/inv_0/op x4in 0.04fF
C1255 cla_1/nand_0/w_0_0# gnd 0.01fF
C1256 cla_0/n nor_1/w_0_0# 0.06fF
C1257 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.06fF
C1258 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/inv_1/w_0_6# 0.03fF
C1259 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.31fF
C1260 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.32fF
C1261 ffo_0/nand_7/a vdd 0.30fF
C1262 vdd ffo_0/nand_1/w_0_0# 0.10fF
C1263 vdd sumffo_2/ffo_0/nand_5/w_0_0# 0.10fF
C1264 vdd sumffo_2/ffo_0/inv_0/op 0.17fF
C1265 gnd cla_2/n 0.22fF
C1266 gnd ffipgarr_0/ffi_0/inv_0/op 0.10fF
C1267 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C1268 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_0/q 0.73fF
C1269 ffipgarr_0/ffipg_1/ffi_1/inv_0/op ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# 0.03fF
C1270 ffipgarr_0/ffipg_0/ffi_0/q nand_5/a 0.02fF
C1271 vdd inv_2/in 0.09fF
C1272 nor_0/a ffipgarr_0/ffipg_0/ffi_1/q 0.22fF
C1273 vdd cla_0/g0 0.50fF
C1274 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/ffi_0/q 0.12fF
C1275 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/a 0.31fF
C1276 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C1277 x3in ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# 0.06fF
C1278 ffipgarr_0/ffipg_1/ffi_1/inv_0/op x2in 0.04fF
C1279 cla_0/inv_0/op cla_0/inv_0/w_0_6# 0.03fF
C1280 inv_6/in nor_4/a 0.04fF
C1281 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/nand_1/a 0.13fF
C1282 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.06fF
C1283 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# sumffo_3/k 0.21fF
C1284 ffipgarr_0/ffipg_0/ffi_1/nand_3/a ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.06fF
C1285 vdd ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# 0.10fF
C1286 vdd sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C1287 vdd ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.17fF
C1288 gnd ffipgarr_0/ffipg_0/ffi_0/nand_0/a_13_n26# 0.01fF
C1289 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.06fF
C1290 nand_2/b cla_0/n 0.05fF
C1291 vdd ffo_0/nand_1/a 0.30fF
C1292 ffipgarr_0/ffipg_1/ffi_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.13fF
C1293 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_0/w_0_0# 0.04fF
C1294 vdd cla_0/nand_0/w_0_0# 0.10fF
C1295 gnd cla_2/nand_0/a_13_n26# 0.01fF
C1296 gnd inv_7/in 0.13fF
C1297 gnd sumffo_3/ffo_0/nand_7/a 0.03fF
C1298 vdd ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# 0.10fF
C1299 ffipgarr_0/ffipg_0/ffi_1/qbar ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.04fF
C1300 cla_1/g0 cla_2/p0 0.32fF
C1301 cla_0/l cla_1/p0 0.02fF
C1302 sumffo_2/ffo_0/nand_3/b vdd 0.39fF
C1303 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.12fF
C1304 ffo_0/inv_0/w_0_6# ffo_0/inv_0/op 0.03fF
C1305 vdd ffo_0/nand_3/b 0.39fF
C1306 ffipgarr_0/ffi_0/nand_1/a clk 0.13fF
C1307 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.30fF
C1308 inv_0/op inv_0/in 0.04fF
C1309 gnd sumffo_1/ffo_0/nand_1/a 0.27fF
C1310 ffipgarr_0/ffipg_0/ffi_1/nand_6/a ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# 0.06fF
C1311 clk nand_5/a 0.11fF
C1312 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.06fF
C1313 clk sumffo_0/ffo_0/nand_5/w_0_0# 0.06fF
C1314 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/op 1.63fF
C1315 clk ffipgarr_0/ffi_0/nand_3/a 0.13fF
C1316 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/q 0.06fF
C1317 vdd ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# 0.10fF
C1318 vdd ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C1319 vdd ffipgarr_0/ffipg_0/ffi_1/nand_7/a 0.34fF
C1320 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C1321 gnd ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# 0.00fF
C1322 nor_0/b ffipgarr_0/ffi_0/nand_6/a 0.00fF
C1323 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C1324 cla_2/l inv_5/w_0_6# 0.29fF
C1325 nand_2/b inv_3/w_0_6# 0.06fF
C1326 sumffo_1/ffo_0/nand_7/w_0_0# vdd 0.10fF
C1327 vdd ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# 0.10fF
C1328 inv_1/w_0_6# inv_1/in 0.10fF
C1329 clk sumffo_0/ffo_0/nand_6/a 0.13fF
C1330 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_1/q 0.73fF
C1331 vdd ffipgarr_0/ffi_0/nand_1/w_0_0# 0.10fF
C1332 ffipgarr_0/ffipg_0/ffi_0/inv_1/op clk 0.07fF
C1333 vdd nor_2/w_0_0# 0.15fF
C1334 nand_0/w_0_0# inv_0/op 0.06fF
C1335 cla_2/p0 cla_2/p1 0.24fF
C1336 y4in ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.01fF
C1337 gnd ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.03fF
C1338 clk ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.07fF
C1339 gnd ffipgarr_0/ffipg_1/ffi_1/nand_1/a 0.14fF
C1340 sumffo_2/ffo_0/nand_6/w_0_0# sumffo_2/sbar 0.04fF
C1341 ffipgarr_0/ffipg_3/ffi_1/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1342 vdd sumffo_3/ffo_0/nand_5/w_0_0# 0.10fF
C1343 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/q 0.06fF
C1344 ffipgarr_0/ffipg_2/ffi_0/nand_3/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.04fF
C1345 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_1/b 0.31fF
C1346 sumffo_1/ffo_0/nand_0/b sumffo_1/ffo_0/d 0.40fF
C1347 gnd cla_1/n 0.08fF
C1348 cla_0/n sumffo_3/k 0.05fF
C1349 clk sumffo_1/ffo_0/nand_5/w_0_0# 0.06fF
C1350 gnd ffipgarr_0/ffipg_3/ffi_1/nand_3/a 0.03fF
C1351 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C1352 cla_1/g0 nand_2/b 1.65fF
C1353 vdd cla_2/g1 0.35fF
C1354 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/op 1.63fF
C1355 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_0/w_0_6# 0.03fF
C1356 inv_2/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1357 sumffo_0/ffo_0/nand_1/b sumffo_0/ffo_0/nand_3/b 0.32fF
C1358 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.04fF
C1359 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_1/ffi_0/q 0.22fF
C1360 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C1361 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.06fF
C1362 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/nand_1/a 0.04fF
C1363 gnd ffo_0/inv_0/op 0.34fF
C1364 clk ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# 0.06fF
C1365 cla_0/l gnd 0.88fF
C1366 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C1367 sumffo_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C1368 ffipgarr_0/ffi_0/nand_4/w_0_0# ffipgarr_0/ffi_0/inv_1/op 0.06fF
C1369 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/qbar 0.32fF
C1370 cla_1/inv_0/op cla_1/nand_0/w_0_0# 0.06fF
C1371 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C1372 sumffo_0/ffo_0/nand_2/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C1373 nor_1/b gnd 0.10fF
C1374 sumffo_1/ffo_0/nand_7/a sumffo_1/ffo_0/nand_5/w_0_0# 0.04fF
C1375 gnd ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.26fF
C1376 nand_2/b cla_1/nor_0/a_13_6# 0.01fF
C1377 vdd ffipgarr_0/ffipg_1/ffi_1/qbar 0.33fF
C1378 sumffo_1/ffo_0/d sumffo_1/xor_0/a_10_10# 0.45fF
C1379 gnd sumffo_1/ffo_0/d 0.37fF
C1380 vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C1381 gnd sumffo_0/ffo_0/nand_1/b 0.26fF
C1382 vdd ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.10fF
C1383 x3in ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# 0.06fF
C1384 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.31fF
C1385 ffipgarr_0/ffipg_0/ffi_0/qbar ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# 0.04fF
C1386 vdd ffipgarr_0/ffi_0/inv_1/op 1.67fF
C1387 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.06fF
C1388 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C1389 vdd cla_0/nor_1/w_0_0# 0.31fF
C1390 nand_2/b inv_3/in 0.13fF
C1391 gnd sumffo_0/ffo_0/nand_7/a 0.03fF
C1392 gnd ffipgarr_0/ffipg_1/ffi_0/nand_0/a_13_n26# 0.01fF
C1393 gnd ffipgarr_0/ffipg_3/ffi_0/nand_1/b 0.26fF
C1394 gnd ffipgarr_0/ffipg_2/ffi_0/nand_1/b 0.26fF
C1395 y1in ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.06fF
C1396 inv_7/op nand_5/a 0.38fF
C1397 cla_2/l inv_7/in 0.13fF
C1398 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C1399 sumffo_3/ffo_0/inv_0/op sumffo_3/ffo_0/nand_0/b 0.32fF
C1400 ffipgarr_0/ffipg_3/ffi_0/qbar ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.00fF
C1401 vdd ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.10fF
C1402 ffipgarr_0/ffipg_1/ffi_1/nand_1/b ffipgarr_0/ffipg_1/ffi_1/inv_1/op 0.45fF
C1403 sumffo_1/sbar sumffo_1/ffo_0/nand_6/w_0_0# 0.04fF
C1404 gnd ffo_0/nand_6/a 0.03fF
C1405 nand_0/w_0_0# nand_2/b 0.04fF
C1406 clk sumffo_3/ffo_0/nand_0/b 0.04fF
C1407 sumffo_3/k ffipgarr_0/ffipg_3/pggen_0/nor_0/a_13_6# 0.01fF
C1408 nand_2/b inv_1/in 0.04fF
C1409 ffo_0/d nor_4/w_0_0# 0.03fF
C1410 vdd sumffo_2/ffo_0/nand_1/b 0.31fF
C1411 vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/a 0.34fF
C1412 vdd ffipgarr_0/ffi_0/inv_1/w_0_6# 0.06fF
C1413 ffipgarr_0/ffipg_2/ffi_1/nand_1/a ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.31fF
C1414 vdd cla_0/inv_0/op 0.17fF
C1415 sumffo_2/ffo_0/nand_6/a sumffo_2/sbar 0.00fF
C1416 sumffo_2/ffo_0/nand_0/w_0_0# sumffo_2/ffo_0/inv_0/op 0.06fF
C1417 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C1418 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C1419 ffo_0/inv_1/w_0_6# ffo_0/nand_0/b 0.03fF
C1420 gnd ffipgarr_0/ffipg_2/ffi_0/nand_7/a 0.03fF
C1421 gnd ffipgarr_0/ffipg_1/ffi_0/nand_6/a 0.03fF
C1422 cla_0/n nor_2/b 0.22fF
C1423 sumffo_2/sbar z3o 0.32fF
C1424 vdd sumffo_0/xor_0/inv_1/op 0.15fF
C1425 vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/a 0.34fF
C1426 vdd cla_1/p0 0.44fF
C1427 ffo_0/inv_0/w_0_6# vdd 0.06fF
C1428 vdd sumffo_1/sbar 0.28fF
C1429 vdd ffipgarr_0/ffi_0/nand_2/w_0_0# 0.10fF
C1430 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_3/w_0_0# 0.04fF
C1431 vdd sumffo_2/ffo_0/nand_1/w_0_0# 0.10fF
C1432 gnd ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.22fF
C1433 ffipgarr_0/ffipg_0/ffi_0/nand_1/a gnd 0.14fF
C1434 cla_0/g0 nand_5/a 0.05fF
C1435 gnd couto 0.52fF
C1436 ffipgarr_0/ffipg_3/ffi_1/nand_6/a ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.13fF
C1437 vdd ffo_0/nand_3/a 0.30fF
C1438 ffipgarr_0/ffi_0/inv_0/op ffipgarr_0/ffi_0/inv_0/w_0_6# 0.03fF
C1439 ffipgarr_0/ffipg_0/ffi_0/q cla_0/g0 1.40fF
C1440 cla_0/l nor_0/a 0.16fF
C1441 vdd cla_1/l 0.27fF
C1442 sumffo_0/ffo_0/nand_3/w_0_0# sumffo_0/ffo_0/nand_3/b 0.06fF
C1443 vdd nor_3/w_0_0# 0.17fF
C1444 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.30fF
C1445 gnd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.17fF
C1446 ffipgarr_0/ffipg_1/ffi_1/nand_6/a ffipgarr_0/ffipg_1/ffi_1/qbar 0.00fF
C1447 ffipgarr_0/ffipg_1/ffi_1/inv_0/op clk 0.32fF
C1448 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# 0.16fF
C1449 sumffo_2/ffo_0/inv_0/op sumffo_2/ffo_0/d 0.04fF
C1450 vdd sumffo_0/ffo_0/d 0.04fF
C1451 vdd ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# 0.11fF
C1452 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.32fF
C1453 inv_4/in nor_2/w_0_0# 0.11fF
C1454 vdd sumffo_1/ffo_0/nand_0/b 0.15fF
C1455 sumffo_1/ffo_0/d sumffo_1/ffo_0/inv_0/w_0_6# 0.06fF
C1456 cla_0/l cla_2/l 0.40fF
C1457 ffo_0/qbar ffo_0/nand_6/a 0.00fF
C1458 cla_2/p1 sumffo_3/k 0.05fF
C1459 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.06fF
C1460 gnd inv_5/in 0.17fF
C1461 nand_2/b ffipgarr_0/ffipg_1/ffi_0/q 0.32fF
C1462 inv_3/w_0_6# nor_2/b 0.03fF
C1463 inv_2/op gnd 0.26fF
C1464 vdd sumffo_0/ffo_0/nand_3/b 0.39fF
C1465 gnd ffipgarr_0/ffipg_2/ffi_1/nand_0/a_13_n26# 0.01fF
C1466 vdd cinin 0.04fF
C1467 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C1468 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/ffi_0/q 0.20fF
C1469 vdd y1in 0.04fF
C1470 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C1471 cla_0/n inv_5/w_0_6# 0.06fF
C1472 gnd sumffo_0/sbar 0.34fF
C1473 gnd ffipgarr_0/ffi_0/nand_7/a 0.03fF
C1474 cla_1/nor_1/w_0_0# cla_2/g0 0.02fF
C1475 cla_1/nand_0/w_0_0# cla_0/n 0.01fF
C1476 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.04fF
C1477 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C1478 vdd ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.10fF
C1479 vdd ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# 0.06fF
C1480 vdd ffipgarr_0/ffipg_1/ffi_0/nand_7/a 0.34fF
C1481 z3o sumffo_2/ffo_0/nand_7/a 0.00fF
C1482 clk sumffo_2/ffo_0/nand_5/w_0_0# 0.06fF
C1483 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.00fF
C1484 sumffo_2/k ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.06fF
C1485 cla_2/g1 cla_2/inv_0/op 0.35fF
C1486 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.04fF
C1487 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C1488 cla_0/g0 clk 0.10fF
C1489 ffo_0/qbar couto 0.32fF
C1490 vdd sumffo_1/xor_0/a_10_10# 0.93fF
C1491 vdd ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# 0.10fF
C1492 gnd ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.03fF
C1493 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C1494 gnd ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.35fF
C1495 vdd gnd 7.04fF
C1496 vdd ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C1497 ffipgarr_0/ffi_0/nand_1/a ffipgarr_0/ffi_0/nand_1/w_0_0# 0.06fF
C1498 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C1499 sumffo_3/sbar sumffo_3/ffo_0/nand_6/a 0.00fF
C1500 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C1501 ffipgarr_0/ffipg_1/ffi_0/nand_1/a ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.31fF
C1502 sumffo_2/k inv_2/op 0.09fF
C1503 sumffo_2/ffo_0/nand_7/w_0_0# vdd 0.10fF
C1504 vdd ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# 0.10fF
C1505 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C1506 clk sumffo_3/ffo_0/inv_1/w_0_6# 0.06fF
C1507 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# 0.06fF
C1508 ffipgarr_0/ffipg_2/ffi_0/inv_1/op ffipgarr_0/ffipg_2/ffi_0/nand_3/b 0.33fF
C1509 clk ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.32fF
C1510 vdd ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# 0.10fF
C1511 sumffo_1/ffo_0/nand_3/b sumffo_1/ffo_0/nand_1/b 0.32fF
C1512 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_2/ffi_1/nand_1/b 0.06fF
C1513 ffipgarr_0/ffipg_2/ffi_0/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op 0.22fF
C1514 ffo_0/nand_0/w_0_0# ffo_0/nand_0/b 0.06fF
C1515 ffipgarr_0/ffipg_3/ffi_0/q ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.31fF
C1516 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/ffi_0/q 0.23fF
C1517 vdd ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# 0.10fF
C1518 sumffo_1/k nand_2/b 0.51fF
C1519 sumffo_1/k ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C1520 inv_3/in nor_2/b 0.04fF
C1521 sumffo_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C1522 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/a 0.30fF
C1523 vdd ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# 0.10fF
C1524 ffo_0/nand_4/w_0_0# ffo_0/nand_6/a 0.04fF
C1525 ffipgarr_0/ffipg_0/ffi_0/nand_1/b ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# 0.06fF
C1526 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# clk 0.06fF
C1527 x1in ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# 0.06fF
C1528 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op gnd 0.17fF
C1529 sumffo_2/ffo_0/nand_3/b clk 0.33fF
C1530 vdd sumffo_2/ffo_0/nand_3/w_0_0# 0.11fF
C1531 sumffo_2/k vdd 0.29fF
C1532 vdd ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C1533 clk ffo_0/nand_3/b 0.33fF
C1534 vdd sumffo_3/ffo_0/nand_4/w_0_0# 0.10fF
C1535 clk ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.13fF
C1536 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.27fF
C1537 sumffo_2/k sumffo_2/xor_0/inv_1/op 0.06fF
C1538 ffipgarr_0/ffipg_2/ffi_1/inv_0/op ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# 0.03fF
C1539 gnd x2in 0.19fF
C1540 cla_2/p0 cla_2/g0 0.15fF
C1541 cla_0/l sumffo_2/ffo_0/nand_3/a 0.15fF
C1542 ffo_0/qbar vdd 0.28fF
C1543 ffo_0/nand_5/w_0_0# ffo_0/nand_1/b 0.06fF
C1544 sumffo_3/k sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C1545 sumffo_3/ffo_0/nand_0/b sumffo_3/ffo_0/inv_1/w_0_6# 0.03fF
C1546 clk ffipgarr_0/ffipg_3/ffi_1/inv_1/op 0.07fF
C1547 ffipgarr_0/ffipg_1/ffi_0/q ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# 0.06fF
C1548 vdd ffipgarr_0/ffipg_0/ffi_0/qbar 0.33fF
C1549 sumffo_3/ffo_0/nand_1/a sumffo_3/ffo_0/nand_3/b 0.00fF
C1550 vdd sumffo_0/ffo_0/inv_0/w_0_6# 0.06fF
C1551 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.04fF
C1552 gnd ffo_0/nand_2/a_13_n26# 0.01fF
C1553 cla_2/l inv_5/in 0.03fF
C1554 gnd ffipgarr_0/ffipg_1/ffi_1/nand_6/a 0.03fF
C1555 ffipgarr_0/ffipg_1/ffi_1/q ffipgarr_0/ffipg_1/ffi_0/q 0.73fF
C1556 vdd ffipgarr_0/ffipg_3/ffi_1/nand_1/b 0.31fF
C1557 ffipgarr_0/ffipg_0/ffi_1/q ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# 0.04fF
C1558 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# clk 0.06fF
C1559 inv_8/w_0_6# inv_8/in 0.10fF
C1560 cla_0/n sumffo_2/ffo_0/nand_4/w_0_0# 0.24fF
C1561 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.06fF
C1562 inv_6/in cla_2/n 0.02fF
C1563 vdd sumffo_1/ffo_0/inv_0/w_0_6# 0.08fF
C1564 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.30fF
C1565 vdd ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# 0.11fF
C1566 vdd nor_0/a 0.29fF
C1567 ffipgarr_0/ffipg_2/ffi_1/nand_7/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.31fF
C1568 sumffo_3/ffo_0/d sumffo_3/xor_0/inv_0/op 0.06fF
C1569 clk sumffo_3/ffo_0/nand_5/w_0_0# 0.06fF
C1570 vdd sumffo_1/ffo_0/nand_3/a 0.30fF
C1571 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/d 0.04fF
C1572 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# sumffo_3/k 0.45fF
C1573 gnd ffipgarr_0/ffipg_2/ffi_0/qbar 0.34fF
C1574 vdd ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# 0.06fF
C1575 vdd ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C1576 cla_0/n cla_1/n 0.09fF
C1577 sumffo_2/ffo_0/d sumffo_2/xor_0/w_n3_4# 0.02fF
C1578 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.06fF
C1579 nor_4/a inv_9/in 0.02fF
C1580 sumffo_1/ffo_0/nand_7/w_0_0# sumffo_1/ffo_0/nand_7/a 0.06fF
C1581 vdd ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# 0.11fF
C1582 vdd ffipgarr_0/ffipg_2/ffi_1/q 1.35fF
C1583 ffipgarr_0/ffipg_1/ffi_0/inv_1/op clk 0.07fF
C1584 vdd cla_2/l 0.40fF
C1585 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/a 0.00fF
C1586 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C1587 vdd ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# 0.06fF
C1588 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op 0.17fF
C1589 gnd ffipgarr_0/ffipg_0/ffi_0/nand_6/a 0.03fF
C1590 gnd ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# 0.01fF
C1591 cla_0/l cla_0/n 0.83fF
C1592 cla_1/p0 nand_5/a 0.00fF
C1593 sumffo_3/ffo_0/d sumffo_3/xor_0/w_n3_4# 0.02fF
C1594 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C1595 sumffo_0/xor_0/inv_1/op nand_5/a 0.22fF
C1596 ffipgarr_0/ffipg_0/ffi_0/inv_0/op ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# 0.03fF
C1597 vdd sumffo_3/ffo_0/nand_1/w_0_0# 0.10fF
C1598 vdd sumffo_2/ffo_0/nand_0/b 0.15fF
C1599 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.04fF
C1600 vdd sumffo_2/ffo_0/inv_1/w_0_6# 0.06fF
C1601 ffipgarr_0/ffi_0/nand_2/w_0_0# ffipgarr_0/ffi_0/nand_3/a 0.04fF
C1602 sumffo_3/ffo_0/nand_1/b sumffo_3/ffo_0/nand_7/a 0.13fF
C1603 sumffo_3/ffo_0/nand_3/a sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C1604 sumffo_0/ffo_0/nand_0/w_0_0# sumffo_0/ffo_0/nand_0/b 0.06fF
C1605 nor_1/b cla_0/n 0.37fF
C1606 ffo_0/nand_4/w_0_0# vdd 0.10fF
C1607 gnd ffipgarr_0/ffipg_3/ffi_1/nand_6/a 0.03fF
C1608 gnd sumffo_0/ffo_0/inv_0/op 0.10fF
C1609 gnd inv_4/in 0.24fF
C1610 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_0/op 0.06fF
C1611 vdd ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# 0.06fF
C1612 ffipgarr_0/ffipg_3/ffi_0/inv_1/op ffipgarr_0/ffipg_3/ffi_0/nand_6/a 0.13fF
C1613 clk ffipgarr_0/ffi_0/inv_1/op 0.10fF
C1614 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.06fF
C1615 sumffo_1/k ffipgarr_0/ffipg_1/ffi_1/q 0.46fF
C1616 vdd cla_1/inv_0/op 0.17fF
C1617 vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.34fF
C1618 gnd cla_2/inv_0/op 0.10fF
C1619 ffipgarr_0/ffipg_2/ffi_0/nand_6/a ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# 0.04fF
C1620 gnd nor_4/b 0.67fF
C1621 ffipgarr_0/ffipg_0/ffi_1/inv_1/op ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.13fF
C1622 ffo_0/nand_1/w_0_0# ffo_0/nand_1/a 0.06fF
C1623 vdd ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# 0.10fF
C1624 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.39fF
C1625 sumffo_3/ffo_0/nand_3/b sumffo_3/ffo_0/nand_3/w_0_0# 0.06fF
C1626 ffipgarr_0/ffipg_3/ffi_1/qbar ffipgarr_0/ffipg_3/ffi_1/q 0.32fF
C1627 cla_0/l inv_3/w_0_6# 0.17fF
C1628 cla_2/g1 cla_2/inv_0/in 0.04fF
C1629 gnd ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C1630 clk sumffo_2/ffo_0/nand_1/b 0.45fF
C1631 ffipgarr_0/ffipg_3/ffi_1/q sumffo_3/k 0.46fF
C1632 clk ffipgarr_0/ffi_0/inv_1/w_0_6# 0.06fF
C1633 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C1634 vdd ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# 0.10fF
C1635 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_3/b 0.04fF
C1636 ffo_0/nand_1/w_0_0# ffo_0/nand_3/b 0.04fF
C1637 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_3/ffi_0/nand_1/a 0.04fF
C1638 vdd ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# 0.11fF
C1639 vdd ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C1640 vdd ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# 0.10fF
C1641 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# ffipgarr_0/ffipg_1/ffi_0/nand_3/a 0.04fF
C1642 ffipgarr_0/ffipg_2/ffi_1/nand_6/a ffipgarr_0/ffipg_2/ffi_1/qbar 0.00fF
C1643 ffipgarr_0/ffipg_0/ffi_0/nand_6/a ffipgarr_0/ffipg_0/ffi_0/qbar 0.00fF
C1644 vdd ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# 0.10fF
C1645 ffipgarr_0/ffipg_3/ffi_0/q sumffo_3/k 0.07fF
C1646 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_3/ffi_0/q 0.23fF
C1647 gnd ffipgarr_0/ffi_0/nand_1/a 0.14fF
C1648 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# ffipgarr_0/ffipg_1/ffi_0/qbar 0.04fF
C1649 vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# 0.06fF
C1650 ffipgarr_0/ffipg_0/ffi_0/inv_1/op y1in 0.01fF
C1651 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C1652 vdd sumffo_1/ffo_0/nand_3/w_0_0# 0.11fF
C1653 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_3/ffi_1/qbar 0.04fF
C1654 ffipgarr_0/ffi_0/nand_2/w_0_0# clk 0.06fF
C1655 vdd ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# 0.10fF
C1656 vdd cla_1/inv_0/in 0.05fF
C1657 ffipgarr_0/ffipg_3/ffi_0/nand_3/b ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# 0.04fF
C1658 ffipgarr_0/ffipg_2/ffi_1/q ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# 0.04fF
C1659 gnd nand_5/a 0.91fF
C1660 cla_2/g0 sumffo_3/k 0.10fF
C1661 cla_2/p1 cla_2/nor_0/w_0_0# 0.06fF
C1662 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# sumffo_3/k 0.02fF
C1663 sumffo_0/ffo_0/nand_1/w_0_0# sumffo_0/ffo_0/nand_3/b 0.04fF
C1664 vdd cla_2/nor_1/w_0_0# 0.31fF
C1665 gnd ffipgarr_0/ffi_0/nand_3/a 0.03fF
C1666 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/inv_0/op 0.06fF
C1667 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# ffipgarr_0/ffipg_1/ffi_1/nand_3/b 0.06fF
C1668 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C1669 ffipgarr_0/ffipg_0/ffi_0/q gnd 2.63fF
C1670 vdd sumffo_2/ffo_0/nand_3/a 0.30fF
C1671 sumffo_0/ffo_0/inv_0/op sumffo_0/ffo_0/inv_0/w_0_6# 0.03fF
C1672 clk ffipgarr_0/ffipg_3/ffi_1/nand_1/a 0.13fF
C1673 vdd ffipgarr_0/ffi_0/inv_0/w_0_6# 0.06fF
C1674 vdd ffipgarr_0/ffipg_0/ffi_1/qbar 0.33fF
C1675 vdd ffipgarr_0/ffipg_0/ffi_0/inv_0/op 0.17fF
C1676 clk sumffo_0/ffo_0/d 0.25fF
C1677 ffo_0/nand_3/b ffo_0/nand_1/a 0.00fF
C1678 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C1679 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C1680 sumffo_1/ffo_0/inv_0/op sumffo_1/ffo_0/nand_0/w_0_0# 0.06fF
C1681 gnd sumffo_0/ffo_0/nand_6/a 0.03fF
C1682 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# ffipgarr_0/ffipg_2/ffi_1/qbar 0.04fF
C1683 ffipgarr_0/ffipg_0/ffi_0/inv_1/op gnd 0.22fF
C1684 sumffo_3/ffo_0/inv_0/w_0_6# vdd 0.06fF
C1685 vdd ffipgarr_0/ffipg_0/ffi_1/nand_6/a 0.34fF
C1686 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_1/b 0.31fF
C1687 ffipgarr_0/ffipg_0/ffi_1/nand_1/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.06fF
C1688 ffo_0/nand_2/w_0_0# ffo_0/nand_0/b 0.06fF
C1689 clk sumffo_1/ffo_0/nand_0/b 0.04fF
C1690 sumffo_1/sbar sumffo_1/ffo_0/nand_7/a 0.31fF
C1691 gnd sumffo_2/ffo_0/d 0.37fF
C1692 gnd ffipgarr_0/ffipg_2/ffi_1/inv_1/op 0.22fF
C1693 clk sumffo_0/ffo_0/nand_3/b 0.33fF
C1694 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# ffipgarr_0/ffipg_3/ffi_1/nand_3/b 0.04fF
C1695 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# ffipgarr_0/ffipg_3/ffi_0/inv_1/op 0.06fF
C1696 clk cinin 0.70fF
C1697 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_2/ffi_0/nand_1/a 0.04fF
C1698 y1in clk 0.70fF
C1699 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# ffipgarr_0/ffipg_0/ffi_0/nand_1/a 0.04fF
C1700 cla_0/n inv_5/in 0.13fF
C1701 inv_2/op cla_0/n 0.70fF
C1702 cla_0/l inv_3/in 0.06fF
C1703 sumffo_2/ffo_0/nand_1/b sumffo_2/ffo_0/nand_1/a 0.31fF
C1704 vdd ffipgarr_0/ffi_0/nand_6/w_0_0# 0.10fF
C1705 sumffo_0/k ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C1706 vdd sumffo_0/ffo_0/nand_0/b 0.15fF
C1707 vdd ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# 0.11fF
C1708 vdd ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# 0.10fF
C1709 gnd sumffo_3/ffo_0/inv_0/op 0.32fF
C1710 ffipgarr_0/ffipg_2/ffi_0/q cla_2/g0 0.13fF
C1711 ffipgarr_0/ffipg_0/ffi_1/nand_1/a ffipgarr_0/ffipg_0/ffi_1/nand_3/b 0.00fF
C1712 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# 0.04fF
C1713 nor_3/b nor_3/w_0_0# 0.06fF
C1714 vdd ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# 0.10fF
C1715 ffipgarr_0/ffipg_1/ffi_1/nand_1/a ffipgarr_0/ffipg_1/ffi_1/nand_1/b 0.31fF
C1716 vdd y2in 0.04fF
C1717 vdd ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# 0.10fF
C1718 clk ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# 0.06fF
C1719 vdd nor_0/w_0_0# 0.15fF
C1720 sumffo_2/ffo_0/nand_1/a sumffo_2/ffo_0/nand_1/w_0_0# 0.06fF
C1721 gnd ffipgarr_0/ffipg_2/ffi_0/nand_6/a 0.03fF
C1722 gnd clk 8.12fF
C1723 cla_0/l inv_1/in 0.08fF
C1724 ffipgarr_0/ffipg_2/ffi_0/nand_1/b ffipgarr_0/ffipg_2/ffi_0/inv_1/op 0.45fF
C1725 vdd ffipgarr_0/ffipg_1/ffi_1/nand_3/a 0.30fF
C1726 ffipgarr_0/ffipg_1/ffi_0/nand_7/a ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# 0.06fF
C1727 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/qbar 0.32fF
C1728 vdd cla_0/n 0.68fF
C1729 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.08fF
C1730 nor_1/b inv_1/in 0.04fF
C1731 ffipgarr_0/ffipg_1/ffi_1/nand_3/a ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# 0.06fF
C1732 nor_0/a nand_5/a 0.26fF
C1733 sumffo_3/ffo_0/nand_2/w_0_0# vdd 0.10fF
C1734 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C1735 gnd z4o 0.52fF
C1736 vdd sumffo_3/ffo_0/nand_0/w_0_0# 0.10fF
C1737 sumffo_1/ffo_0/nand_6/a sumffo_1/ffo_0/nand_4/w_0_0# 0.04fF
C1738 ffipgarr_0/ffipg_0/ffi_0/q nor_0/a 0.14fF
C1739 gnd sumffo_1/ffo_0/nand_7/a 0.03fF
C1740 ffipgarr_0/ffipg_2/ffi_1/nand_3/b ffipgarr_0/ffipg_2/ffi_1/nand_3/a 0.31fF
C1741 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C1742 inv_1/w_0_6# nand_2/b 0.01fF
C1743 vdd nor_4/w_0_0# 0.15fF
C1744 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# 0.16fF
C1745 vdd ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# 0.10fF
C1746 sumffo_0/k nor_0/b 0.09fF
C1747 sumffo_2/ffo_0/nand_5/w_0_0# sumffo_2/ffo_0/nand_1/b 0.06fF
C1748 ffipgarr_0/ffipg_2/ffi_1/nand_1/a clk 0.13fF
C1749 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# clk 0.06fF
C1750 nor_3/b gnd 0.10fF
C1751 gnd sumffo_3/ffo_0/nand_0/b 0.38fF
C1752 vdd sumffo_0/ffo_0/inv_1/w_0_6# 0.06fF
C1753 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# ffipgarr_0/ffipg_0/ffi_1/inv_1/op 0.06fF
C1754 vdd inv_3/w_0_6# 0.15fF
C1755 sumffo_3/xor_0/inv_0/op inv_4/op 0.20fF
C1756 clk sumffo_3/ffo_0/nand_4/w_0_0# 0.06fF
C1757 ffo_0/d inv_9/in 0.04fF
C1758 sumffo_3/xor_0/a_10_10# sumffo_3/ffo_0/d 0.45fF
C1759 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/nand_0/w_0_0# 0.06fF
C1760 sumffo_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C1761 gnd cla_2/inv_0/in 0.35fF
C1762 gnd ffipgarr_0/ffipg_3/ffi_0/nand_3/b 0.35fF
C1763 sumffo_3/k sumffo_3/xor_0/inv_0/op 0.27fF
C1764 gnd sumffo_2/ffo_0/nand_1/a 0.06fF
C1765 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# ffipgarr_0/ffipg_0/ffi_1/q 0.06fF
C1766 cla_0/g0 cla_1/p0 0.33fF
C1767 nand_2/b cla_2/p0 0.00fF
C1768 vdd x3in 0.04fF
C1769 vdd y3in 0.04fF
C1770 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op 0.03fF
C1771 ffipgarr_0/ffi_0/nand_3/b ffipgarr_0/ffi_0/nand_3/w_0_0# 0.06fF
C1772 cla_1/nand_0/w_0_0# cla_2/g0 0.06fF
C1773 sumffo_3/xor_0/w_n3_4# inv_4/op 0.06fF
C1774 sumffo_2/ffo_0/nand_6/a sumffo_2/ffo_0/nand_6/w_0_0# 0.06fF
C1775 nor_0/a clk 0.13fF
C1776 vdd sumffo_2/ffo_0/inv_0/w_0_6# 0.06fF
C1777 clk ffipgarr_0/ffipg_2/ffi_0/nand_3/a 0.13fF
C1778 vdd ffipgarr_0/ffipg_1/ffi_0/nand_1/b 0.31fF
C1779 vdd cla_1/g0 0.49fF
C1780 cla_0/inv_0/op cla_0/nand_0/w_0_0# 0.06fF
C1781 vdd inv_6/in 0.09fF
C1782 vdd sumffo_3/ffo_0/nand_1/b 0.31fF
C1783 vdd ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# 0.10fF
C1784 ffipgarr_0/ffipg_0/ffi_0/q ffipgarr_0/ffipg_0/ffi_0/nand_7/a 0.00fF
C1785 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C1786 gnd ffipgarr_0/ffipg_1/ffi_1/inv_0/op 0.10fF
C1787 inv_7/op gnd 0.16fF
C1788 sumffo_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C1789 sumffo_2/ffo_0/nand_6/w_0_0# z3o 0.06fF
C1790 sumffo_2/ffo_0/nand_0/b sumffo_2/ffo_0/d 0.40fF
C1791 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# clk 0.06fF
C1792 ffipgarr_0/ffipg_0/ffi_1/nand_3/b ffipgarr_0/ffipg_0/ffi_1/nand_3/a 0.31fF
C1793 sumffo_2/ffo_0/nand_3/b sumffo_2/ffo_0/nand_1/b 0.32fF
C1794 cla_0/l sumffo_2/ffo_0/nand_2/w_0_0# 0.17fF
C1795 ffipgarr_0/ffipg_0/ffi_1/q nor_0/b 1.27fF
C1796 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C1797 ffipgarr_0/ffipg_3/ffi_1/nand_3/b ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# 0.06fF
C1798 ffipgarr_0/ffipg_3/ffi_0/nand_1/b ffipgarr_0/ffipg_3/ffi_0/nand_7/a 0.13fF
C1799 clk ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# 0.06fF
C1800 ffipgarr_0/ffipg_1/ffi_0/nand_3/b ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# 0.06fF
C1801 vdd ffipgarr_0/ffipg_0/ffi_1/inv_0/op 0.17fF
C1802 inv_9/in Gnd 0.23fF
C1803 nor_4/w_0_0# Gnd 1.81fF
C1804 nor_4/b Gnd 1.06fF
C1805 inv_8/in Gnd 0.22fF
C1806 inv_8/w_0_6# Gnd 1.40fF
C1807 inv_7/in Gnd 0.22fF
C1808 inv_7/w_0_6# Gnd 1.40fF
C1809 nor_4/a Gnd 0.27fF
C1810 inv_5/in Gnd 0.22fF
C1811 inv_5/w_0_6# Gnd 1.40fF
C1812 nor_3/b Gnd 0.92fF
C1813 cla_2/n Gnd 0.32fF
C1814 inv_6/in Gnd 0.23fF
C1815 nor_3/w_0_0# Gnd 1.81fF
C1816 nor_2/b Gnd 0.92fF
C1817 cla_1/n Gnd 0.20fF
C1818 inv_4/in Gnd 0.23fF
C1819 nor_2/w_0_0# Gnd 1.81fF
C1820 inv_3/in Gnd 0.22fF
C1821 inv_3/w_0_6# Gnd 1.40fF
C1822 inv_2/op Gnd 1.94fF
C1823 inv_2/in Gnd 0.23fF
C1824 nor_1/w_0_0# Gnd 1.81fF
C1825 nor_1/b Gnd 0.85fF
C1826 inv_1/in Gnd 0.22fF
C1827 inv_1/w_0_6# Gnd 1.40fF
C1828 inv_0/in Gnd 0.23fF
C1829 nor_0/w_0_0# Gnd 1.81fF
C1830 ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1831 ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1832 ffo_0/nand_7/a Gnd 0.30fF
C1833 ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1834 ffo_0/qbar Gnd 0.42fF
C1835 ffo_0/nand_6/a Gnd 0.30fF
C1836 ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1837 ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1838 ffo_0/nand_3/b Gnd 0.43fF
C1839 ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1840 ffo_0/nand_3/a Gnd 0.30fF
C1841 ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1842 ffo_0/nand_0/b Gnd 0.63fF
C1843 ffo_0/d Gnd 0.60fF
C1844 ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1845 ffo_0/inv_0/op Gnd 0.26fF
C1846 ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1847 ffo_0/nand_1/a Gnd 0.30fF
C1848 ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1849 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C1850 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C1851 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C1852 inv_4/op Gnd 1.54fF
C1853 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1854 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C1855 sumffo_3/k Gnd 3.28fF
C1856 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1857 sumffo_3/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1858 sumffo_3/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1859 sumffo_3/ffo_0/nand_7/a Gnd 0.30fF
C1860 sumffo_3/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1861 sumffo_3/sbar Gnd 0.43fF
C1862 sumffo_3/ffo_0/nand_6/a Gnd 0.30fF
C1863 sumffo_3/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1864 sumffo_3/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1865 sumffo_3/ffo_0/nand_3/b Gnd 0.43fF
C1866 sumffo_3/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1867 sumffo_3/ffo_0/nand_3/a Gnd 0.30fF
C1868 sumffo_3/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1869 sumffo_3/ffo_0/nand_0/b Gnd 0.63fF
C1870 sumffo_3/ffo_0/d Gnd 0.64fF
C1871 sumffo_3/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1872 sumffo_3/ffo_0/inv_0/op Gnd 0.26fF
C1873 sumffo_3/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1874 sumffo_3/ffo_0/nand_1/a Gnd 0.30fF
C1875 sumffo_3/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1876 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C1877 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C1878 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C1879 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1880 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C1881 sumffo_1/k Gnd 2.61fF
C1882 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1883 sumffo_1/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1884 sumffo_1/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1885 sumffo_1/ffo_0/nand_7/a Gnd 0.30fF
C1886 sumffo_1/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1887 sumffo_1/sbar Gnd 0.43fF
C1888 sumffo_1/ffo_0/nand_6/a Gnd 0.30fF
C1889 sumffo_1/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1890 sumffo_1/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1891 sumffo_1/ffo_0/nand_3/b Gnd 0.43fF
C1892 sumffo_1/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1893 sumffo_1/ffo_0/nand_3/a Gnd 0.30fF
C1894 sumffo_1/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1895 sumffo_1/ffo_0/nand_0/b Gnd 0.63fF
C1896 sumffo_1/ffo_0/d Gnd 0.64fF
C1897 sumffo_1/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1898 sumffo_1/ffo_0/inv_0/op Gnd 0.26fF
C1899 sumffo_1/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1900 sumffo_1/ffo_0/nand_1/a Gnd 0.30fF
C1901 sumffo_1/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1902 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C1903 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C1904 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C1905 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1906 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C1907 sumffo_2/k Gnd 1.72fF
C1908 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1909 sumffo_2/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1910 sumffo_2/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1911 gnd Gnd 46.05fF
C1912 sumffo_2/ffo_0/nand_7/a Gnd 0.30fF
C1913 sumffo_2/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1914 sumffo_2/sbar Gnd 0.43fF
C1915 vdd Gnd 27.16fF
C1916 sumffo_2/ffo_0/nand_6/a Gnd 0.30fF
C1917 sumffo_2/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1918 sumffo_2/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1919 sumffo_2/ffo_0/nand_3/b Gnd 0.43fF
C1920 sumffo_2/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1921 sumffo_2/ffo_0/nand_3/a Gnd 0.30fF
C1922 sumffo_2/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1923 sumffo_2/ffo_0/nand_0/b Gnd 0.63fF
C1924 sumffo_2/ffo_0/d Gnd 0.64fF
C1925 sumffo_2/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1926 sumffo_2/ffo_0/inv_0/op Gnd 0.26fF
C1927 sumffo_2/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1928 sumffo_2/ffo_0/nand_1/a Gnd 0.30fF
C1929 sumffo_2/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1930 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C1931 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C1932 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C1933 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C1934 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C1935 sumffo_0/k Gnd 3.08fF
C1936 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C1937 sumffo_0/ffo_0/inv_1/w_0_6# Gnd 0.58fF
C1938 sumffo_0/ffo_0/inv_0/w_0_6# Gnd 0.58fF
C1939 sumffo_0/ffo_0/nand_7/a Gnd 0.30fF
C1940 sumffo_0/ffo_0/nand_7/w_0_0# Gnd 0.82fF
C1941 sumffo_0/sbar Gnd 0.43fF
C1942 sumffo_0/ffo_0/nand_6/a Gnd 0.30fF
C1943 sumffo_0/ffo_0/nand_6/w_0_0# Gnd 0.82fF
C1944 sumffo_0/ffo_0/nand_5/w_0_0# Gnd 0.82fF
C1945 sumffo_0/ffo_0/nand_3/b Gnd 0.43fF
C1946 sumffo_0/ffo_0/nand_4/w_0_0# Gnd 0.82fF
C1947 sumffo_0/ffo_0/nand_3/a Gnd 0.30fF
C1948 sumffo_0/ffo_0/nand_3/w_0_0# Gnd 0.82fF
C1949 sumffo_0/ffo_0/nand_0/b Gnd 0.63fF
C1950 sumffo_0/ffo_0/d Gnd 0.64fF
C1951 sumffo_0/ffo_0/nand_2/w_0_0# Gnd 0.82fF
C1952 sumffo_0/ffo_0/inv_0/op Gnd 0.26fF
C1953 sumffo_0/ffo_0/nand_0/w_0_0# Gnd 0.82fF
C1954 sumffo_0/ffo_0/nand_1/a Gnd 0.30fF
C1955 sumffo_0/ffo_0/nand_1/w_0_0# Gnd 0.82fF
C1956 cla_2/p1 Gnd 1.08fF
C1957 cla_2/nor_1/w_0_0# Gnd 1.23fF
C1958 cla_2/nor_0/w_0_0# Gnd 1.23fF
C1959 cla_2/inv_0/in Gnd 0.27fF
C1960 cla_2/inv_0/w_0_6# Gnd 0.58fF
C1961 cla_2/g1 Gnd 0.58fF
C1962 cla_2/inv_0/op Gnd 0.26fF
C1963 cla_2/nand_0/w_0_0# Gnd 0.82fF
C1964 ffipgarr_0/ffipg_3/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C1965 ffipgarr_0/ffipg_3/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C1966 ffipgarr_0/ffipg_3/ffi_1/nand_7/a Gnd 0.30fF
C1967 ffipgarr_0/ffipg_3/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C1968 ffipgarr_0/ffipg_3/ffi_1/qbar Gnd 0.42fF
C1969 ffipgarr_0/ffipg_3/ffi_1/nand_6/a Gnd 0.30fF
C1970 ffipgarr_0/ffipg_3/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C1971 ffipgarr_0/ffipg_3/ffi_1/inv_1/op Gnd 0.89fF
C1972 ffipgarr_0/ffipg_3/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C1973 ffipgarr_0/ffipg_3/ffi_1/nand_3/b Gnd 0.43fF
C1974 ffipgarr_0/ffipg_3/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C1975 ffipgarr_0/ffipg_3/ffi_1/nand_3/a Gnd 0.30fF
C1976 ffipgarr_0/ffipg_3/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C1977 x4in Gnd 0.52fF
C1978 ffipgarr_0/ffipg_3/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C1979 ffipgarr_0/ffipg_3/ffi_1/inv_0/op Gnd 0.26fF
C1980 ffipgarr_0/ffipg_3/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C1981 ffipgarr_0/ffipg_3/ffi_1/nand_1/a Gnd 0.30fF
C1982 ffipgarr_0/ffipg_3/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C1983 ffipgarr_0/ffipg_3/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C1984 ffipgarr_0/ffipg_3/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C1985 ffipgarr_0/ffipg_3/ffi_0/nand_7/a Gnd 0.30fF
C1986 ffipgarr_0/ffipg_3/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C1987 ffipgarr_0/ffipg_3/ffi_0/qbar Gnd 0.42fF
C1988 ffipgarr_0/ffipg_3/ffi_0/nand_6/a Gnd 0.30fF
C1989 ffipgarr_0/ffipg_3/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C1990 ffipgarr_0/ffipg_3/ffi_0/inv_1/op Gnd 0.89fF
C1991 ffipgarr_0/ffipg_3/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C1992 ffipgarr_0/ffipg_3/ffi_0/nand_3/b Gnd 0.43fF
C1993 ffipgarr_0/ffipg_3/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C1994 ffipgarr_0/ffipg_3/ffi_0/nand_3/a Gnd 0.30fF
C1995 ffipgarr_0/ffipg_3/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C1996 y4in Gnd 0.52fF
C1997 ffipgarr_0/ffipg_3/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C1998 ffipgarr_0/ffipg_3/ffi_0/inv_0/op Gnd 0.26fF
C1999 ffipgarr_0/ffipg_3/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2000 ffipgarr_0/ffipg_3/ffi_0/nand_1/a Gnd 0.30fF
C2001 ffipgarr_0/ffipg_3/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2002 ffipgarr_0/ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2003 ffipgarr_0/ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2004 ffipgarr_0/ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2005 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2006 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2007 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2008 ffipgarr_0/ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2009 ffipgarr_0/ffipg_3/ffi_0/q Gnd 2.68fF
C2010 ffipgarr_0/ffipg_3/ffi_1/q Gnd 2.93fF
C2011 ffipgarr_0/ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2012 ffipgarr_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2013 ffipgarr_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2014 ffipgarr_0/ffi_0/nand_7/a Gnd 0.30fF
C2015 ffipgarr_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2016 nor_0/b Gnd 1.09fF
C2017 ffipgarr_0/ffi_0/nand_6/a Gnd 0.30fF
C2018 ffipgarr_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2019 ffipgarr_0/ffi_0/inv_1/op Gnd 0.89fF
C2020 ffipgarr_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2021 ffipgarr_0/ffi_0/nand_3/b Gnd 0.43fF
C2022 ffipgarr_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2023 ffipgarr_0/ffi_0/nand_3/a Gnd 0.30fF
C2024 ffipgarr_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2025 clk Gnd 17.25fF
C2026 cinin Gnd 0.52fF
C2027 ffipgarr_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2028 ffipgarr_0/ffi_0/inv_0/op Gnd 0.26fF
C2029 ffipgarr_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2030 ffipgarr_0/ffi_0/nand_1/a Gnd 0.30fF
C2031 ffipgarr_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2032 ffipgarr_0/ffipg_2/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2033 ffipgarr_0/ffipg_2/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2034 ffipgarr_0/ffipg_2/ffi_1/nand_7/a Gnd 0.30fF
C2035 ffipgarr_0/ffipg_2/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2036 ffipgarr_0/ffipg_2/ffi_1/qbar Gnd 0.42fF
C2037 ffipgarr_0/ffipg_2/ffi_1/nand_6/a Gnd 0.30fF
C2038 ffipgarr_0/ffipg_2/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2039 ffipgarr_0/ffipg_2/ffi_1/inv_1/op Gnd 0.89fF
C2040 ffipgarr_0/ffipg_2/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2041 ffipgarr_0/ffipg_2/ffi_1/nand_3/b Gnd 0.43fF
C2042 ffipgarr_0/ffipg_2/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2043 ffipgarr_0/ffipg_2/ffi_1/nand_3/a Gnd 0.30fF
C2044 ffipgarr_0/ffipg_2/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2045 x3in Gnd 0.52fF
C2046 ffipgarr_0/ffipg_2/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2047 ffipgarr_0/ffipg_2/ffi_1/inv_0/op Gnd 0.26fF
C2048 ffipgarr_0/ffipg_2/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2049 ffipgarr_0/ffipg_2/ffi_1/nand_1/a Gnd 0.30fF
C2050 ffipgarr_0/ffipg_2/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2051 ffipgarr_0/ffipg_2/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2052 ffipgarr_0/ffipg_2/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2053 ffipgarr_0/ffipg_2/ffi_0/nand_7/a Gnd 0.30fF
C2054 ffipgarr_0/ffipg_2/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2055 ffipgarr_0/ffipg_2/ffi_0/qbar Gnd 0.42fF
C2056 ffipgarr_0/ffipg_2/ffi_0/nand_6/a Gnd 0.30fF
C2057 ffipgarr_0/ffipg_2/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2058 ffipgarr_0/ffipg_2/ffi_0/inv_1/op Gnd 0.89fF
C2059 ffipgarr_0/ffipg_2/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2060 ffipgarr_0/ffipg_2/ffi_0/nand_3/b Gnd 0.43fF
C2061 ffipgarr_0/ffipg_2/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2062 ffipgarr_0/ffipg_2/ffi_0/nand_3/a Gnd 0.30fF
C2063 ffipgarr_0/ffipg_2/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2064 y3in Gnd 0.52fF
C2065 ffipgarr_0/ffipg_2/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2066 ffipgarr_0/ffipg_2/ffi_0/inv_0/op Gnd 0.26fF
C2067 ffipgarr_0/ffipg_2/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2068 ffipgarr_0/ffipg_2/ffi_0/nand_1/a Gnd 0.30fF
C2069 ffipgarr_0/ffipg_2/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2070 ffipgarr_0/ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2071 ffipgarr_0/ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2072 ffipgarr_0/ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2073 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2074 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2075 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2076 ffipgarr_0/ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2077 ffipgarr_0/ffipg_2/ffi_0/q Gnd 2.68fF
C2078 ffipgarr_0/ffipg_2/ffi_1/q Gnd 2.93fF
C2079 ffipgarr_0/ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2080 ffipgarr_0/ffipg_1/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2081 ffipgarr_0/ffipg_1/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2082 ffipgarr_0/ffipg_1/ffi_1/nand_7/a Gnd 0.30fF
C2083 ffipgarr_0/ffipg_1/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2084 ffipgarr_0/ffipg_1/ffi_1/qbar Gnd 0.42fF
C2085 ffipgarr_0/ffipg_1/ffi_1/nand_6/a Gnd 0.30fF
C2086 ffipgarr_0/ffipg_1/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2087 ffipgarr_0/ffipg_1/ffi_1/inv_1/op Gnd 0.89fF
C2088 ffipgarr_0/ffipg_1/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2089 ffipgarr_0/ffipg_1/ffi_1/nand_3/b Gnd 0.43fF
C2090 ffipgarr_0/ffipg_1/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2091 ffipgarr_0/ffipg_1/ffi_1/nand_3/a Gnd 0.30fF
C2092 ffipgarr_0/ffipg_1/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2093 x2in Gnd 0.52fF
C2094 ffipgarr_0/ffipg_1/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2095 ffipgarr_0/ffipg_1/ffi_1/inv_0/op Gnd 0.26fF
C2096 ffipgarr_0/ffipg_1/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2097 ffipgarr_0/ffipg_1/ffi_1/nand_1/a Gnd 0.30fF
C2098 ffipgarr_0/ffipg_1/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2099 ffipgarr_0/ffipg_1/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2100 ffipgarr_0/ffipg_1/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2101 ffipgarr_0/ffipg_1/ffi_0/nand_7/a Gnd 0.30fF
C2102 ffipgarr_0/ffipg_1/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2103 ffipgarr_0/ffipg_1/ffi_0/qbar Gnd 0.42fF
C2104 ffipgarr_0/ffipg_1/ffi_0/nand_6/a Gnd 0.30fF
C2105 ffipgarr_0/ffipg_1/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2106 ffipgarr_0/ffipg_1/ffi_0/inv_1/op Gnd 0.89fF
C2107 ffipgarr_0/ffipg_1/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2108 ffipgarr_0/ffipg_1/ffi_0/nand_3/b Gnd 0.43fF
C2109 ffipgarr_0/ffipg_1/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2110 ffipgarr_0/ffipg_1/ffi_0/nand_3/a Gnd 0.30fF
C2111 ffipgarr_0/ffipg_1/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2112 y2in Gnd 0.43fF
C2113 ffipgarr_0/ffipg_1/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2114 ffipgarr_0/ffipg_1/ffi_0/inv_0/op Gnd 0.26fF
C2115 ffipgarr_0/ffipg_1/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2116 ffipgarr_0/ffipg_1/ffi_0/nand_1/a Gnd 0.30fF
C2117 ffipgarr_0/ffipg_1/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2118 ffipgarr_0/ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2119 ffipgarr_0/ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2120 ffipgarr_0/ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2121 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2122 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2123 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2124 ffipgarr_0/ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2125 ffipgarr_0/ffipg_1/ffi_0/q Gnd 2.68fF
C2126 ffipgarr_0/ffipg_1/ffi_1/q Gnd 2.93fF
C2127 ffipgarr_0/ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2128 ffipgarr_0/ffipg_0/ffi_1/inv_1/w_0_6# Gnd 0.58fF
C2129 ffipgarr_0/ffipg_0/ffi_1/inv_0/w_0_6# Gnd 0.58fF
C2130 ffipgarr_0/ffipg_0/ffi_1/nand_7/a Gnd 0.30fF
C2131 ffipgarr_0/ffipg_0/ffi_1/nand_7/w_0_0# Gnd 0.82fF
C2132 ffipgarr_0/ffipg_0/ffi_1/qbar Gnd 0.42fF
C2133 ffipgarr_0/ffipg_0/ffi_1/nand_6/a Gnd 0.30fF
C2134 ffipgarr_0/ffipg_0/ffi_1/nand_6/w_0_0# Gnd 0.82fF
C2135 ffipgarr_0/ffipg_0/ffi_1/inv_1/op Gnd 0.89fF
C2136 ffipgarr_0/ffipg_0/ffi_1/nand_5/w_0_0# Gnd 0.82fF
C2137 ffipgarr_0/ffipg_0/ffi_1/nand_3/b Gnd 0.43fF
C2138 ffipgarr_0/ffipg_0/ffi_1/nand_4/w_0_0# Gnd 0.82fF
C2139 ffipgarr_0/ffipg_0/ffi_1/nand_3/a Gnd 0.30fF
C2140 ffipgarr_0/ffipg_0/ffi_1/nand_3/w_0_0# Gnd 0.82fF
C2141 x1in Gnd 0.42fF
C2142 ffipgarr_0/ffipg_0/ffi_1/nand_2/w_0_0# Gnd 0.82fF
C2143 ffipgarr_0/ffipg_0/ffi_1/inv_0/op Gnd 0.26fF
C2144 ffipgarr_0/ffipg_0/ffi_1/nand_0/w_0_0# Gnd 0.82fF
C2145 ffipgarr_0/ffipg_0/ffi_1/nand_1/a Gnd 0.30fF
C2146 ffipgarr_0/ffipg_0/ffi_1/nand_1/w_0_0# Gnd 0.82fF
C2147 ffipgarr_0/ffipg_0/ffi_0/inv_1/w_0_6# Gnd 0.58fF
C2148 ffipgarr_0/ffipg_0/ffi_0/inv_0/w_0_6# Gnd 0.58fF
C2149 ffipgarr_0/ffipg_0/ffi_0/nand_7/a Gnd 0.30fF
C2150 ffipgarr_0/ffipg_0/ffi_0/nand_7/w_0_0# Gnd 0.82fF
C2151 ffipgarr_0/ffipg_0/ffi_0/qbar Gnd 0.42fF
C2152 ffipgarr_0/ffipg_0/ffi_0/nand_6/a Gnd 0.30fF
C2153 ffipgarr_0/ffipg_0/ffi_0/nand_6/w_0_0# Gnd 0.82fF
C2154 ffipgarr_0/ffipg_0/ffi_0/inv_1/op Gnd 0.89fF
C2155 ffipgarr_0/ffipg_0/ffi_0/nand_5/w_0_0# Gnd 0.82fF
C2156 ffipgarr_0/ffipg_0/ffi_0/nand_3/b Gnd 0.43fF
C2157 ffipgarr_0/ffipg_0/ffi_0/nand_4/w_0_0# Gnd 0.82fF
C2158 ffipgarr_0/ffipg_0/ffi_0/nand_3/a Gnd 0.30fF
C2159 ffipgarr_0/ffipg_0/ffi_0/nand_3/w_0_0# Gnd 0.82fF
C2160 y1in Gnd 0.52fF
C2161 ffipgarr_0/ffipg_0/ffi_0/nand_2/w_0_0# Gnd 0.82fF
C2162 ffipgarr_0/ffipg_0/ffi_0/inv_0/op Gnd 0.26fF
C2163 ffipgarr_0/ffipg_0/ffi_0/nand_0/w_0_0# Gnd 0.82fF
C2164 ffipgarr_0/ffipg_0/ffi_0/nand_1/a Gnd 0.30fF
C2165 ffipgarr_0/ffipg_0/ffi_0/nand_1/w_0_0# Gnd 0.82fF
C2166 ffipgarr_0/ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C2167 ffipgarr_0/ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C2168 ffipgarr_0/ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C2169 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C2170 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C2171 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C2172 ffipgarr_0/ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C2173 ffipgarr_0/ffipg_0/ffi_0/q Gnd 2.68fF
C2174 ffipgarr_0/ffipg_0/ffi_1/q Gnd 2.93fF
C2175 ffipgarr_0/ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C2176 cla_1/nor_1/w_0_0# Gnd 1.23fF
C2177 cla_1/l Gnd 0.31fF
C2178 cla_1/nor_0/w_0_0# Gnd 1.23fF
C2179 cla_1/inv_0/in Gnd 0.27fF
C2180 cla_1/inv_0/w_0_6# Gnd 0.58fF
C2181 cla_1/inv_0/op Gnd 0.26fF
C2182 cla_1/nand_0/w_0_0# Gnd 0.82fF
C2183 inv_7/op Gnd 0.30fF
C2184 cla_0/nor_1/w_0_0# Gnd 1.23fF
C2185 cla_0/l Gnd 7.05fF
C2186 cla_0/nor_0/w_0_0# Gnd 1.23fF
C2187 cla_0/inv_0/in Gnd 0.27fF
C2188 cla_0/inv_0/w_0_6# Gnd 0.58fF
C2189 cla_1/g0 Gnd 2.32fF
C2190 cla_0/inv_0/op Gnd 0.26fF
C2191 cla_0/nand_0/w_0_0# Gnd 0.82fF
C2192 cla_2/l Gnd 1.05fF
C2193 nand_2/b Gnd 0.27fF
C2194 inv_0/op Gnd 0.26fF
C2195 nand_0/w_0_0# Gnd 0.82fF
