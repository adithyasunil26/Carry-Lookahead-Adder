magic
tech scmos
timestamp 1618763462
<< metal1 >>
rect -17 1666 82 1669
rect 87 1666 523 1669
rect 528 1666 743 1669
rect -17 1659 -15 1662
rect -10 1659 740 1662
rect 737 1591 740 1659
rect 965 1592 969 1595
rect 601 1584 615 1587
rect 742 1586 744 1589
rect 601 1560 604 1584
rect 223 1555 599 1558
rect -17 1552 2 1555
rect -17 1480 -2 1483
rect 472 1413 475 1529
rect 507 1487 510 1555
rect 531 1530 615 1533
rect 507 1484 557 1487
rect 513 1395 516 1484
rect 553 1433 558 1436
rect 555 1423 558 1433
rect 611 1420 617 1423
rect 652 1406 654 1409
rect 994 1398 996 1401
rect 513 1392 519 1395
rect 611 1390 612 1393
rect 617 1390 642 1393
rect 767 1392 771 1395
rect 472 1386 501 1389
rect 506 1386 519 1389
rect 550 1367 553 1378
rect 472 1360 494 1363
rect 499 1360 565 1363
rect 574 1361 577 1375
rect 611 1361 620 1364
rect 634 1336 642 1339
rect -17 1273 -2 1276
rect 634 1275 637 1336
rect 472 1272 637 1275
rect -17 1196 -2 1199
rect 472 1129 475 1272
rect 613 1158 616 1169
rect 576 1142 579 1145
rect 572 1136 579 1139
rect 637 1137 640 1140
rect 508 1126 509 1129
rect 572 1126 575 1136
rect 568 1123 575 1126
rect 641 1111 648 1114
rect 637 1108 644 1111
rect 611 1107 637 1108
rect 472 1102 487 1105
rect 492 1102 507 1105
rect 682 1101 685 1114
rect 469 1068 472 1076
rect 501 1074 507 1077
rect 625 1069 628 1074
rect 644 1070 648 1073
rect 706 1069 714 1072
rect 469 1065 476 1068
rect 481 1065 507 1068
rect 630 1064 648 1067
rect 627 1045 648 1048
rect 682 1045 685 1053
rect 694 1015 714 1018
rect 694 1001 697 1015
rect 840 1013 843 1016
rect 1066 1007 1068 1010
rect 472 998 697 1001
rect -17 989 -2 992
rect -17 916 -2 919
rect 472 849 475 998
rect 554 886 576 889
rect 609 878 612 889
rect 568 862 575 865
rect 570 856 575 859
rect 632 857 635 860
rect 494 846 507 849
rect 570 846 573 856
rect 568 843 573 846
rect 641 831 647 834
rect 632 828 644 831
rect 609 827 633 828
rect 472 822 499 825
rect 504 822 507 825
rect 681 821 684 834
rect 469 788 472 796
rect 480 794 507 797
rect 469 785 479 788
rect 484 785 507 788
rect 625 787 628 794
rect 641 790 647 793
rect 705 789 711 792
rect 625 784 647 787
rect 627 765 647 768
rect 681 765 684 773
rect 695 735 711 738
rect 695 716 698 735
rect 837 733 840 736
rect 1063 727 1065 730
rect 472 713 698 716
rect -17 709 -2 712
rect -17 632 -2 635
rect 472 565 475 713
rect 631 606 655 609
rect 607 594 610 605
rect 631 589 634 606
rect 685 596 688 609
rect 715 596 718 610
rect 752 597 755 610
rect 709 593 718 596
rect 648 582 651 585
rect 568 578 573 581
rect 645 578 651 579
rect 567 572 573 575
rect 648 576 651 578
rect 709 577 718 580
rect 567 562 570 572
rect 1008 567 1010 570
rect 565 559 570 562
rect -24 548 -22 551
rect 709 548 718 551
rect 752 548 755 549
rect 685 547 688 548
rect 631 544 638 547
rect 607 543 631 544
rect 472 538 504 541
rect 672 534 675 547
rect 696 531 705 534
rect 739 521 742 534
rect 469 504 472 512
rect 484 510 504 513
rect 469 501 504 504
rect 622 500 625 510
rect 782 508 787 511
rect 634 503 638 506
rect 696 502 702 505
rect 622 497 638 500
rect 699 493 702 502
rect 699 490 705 493
rect 782 492 785 508
rect 763 489 785 492
rect -17 425 -2 428
rect -2 387 58 390
rect 607 390 610 481
rect 621 478 638 481
rect 672 478 675 486
rect 693 468 696 486
rect 693 465 705 468
rect 739 465 742 473
rect 63 387 809 390
<< m2contact >>
rect 472 1529 477 1534
rect 526 1530 531 1535
rect 557 1482 562 1487
rect 647 1405 652 1410
rect 612 1389 617 1394
rect 501 1384 506 1389
rect 575 1383 580 1388
rect 494 1359 499 1364
rect 565 1360 570 1365
rect 620 1361 625 1366
rect 571 1142 576 1147
rect 640 1137 645 1142
rect 503 1126 508 1131
rect 487 1100 492 1105
rect 496 1074 501 1079
rect 639 1070 644 1075
rect 476 1064 481 1069
rect 625 1064 630 1069
rect 563 862 568 867
rect 489 846 494 851
rect 635 855 640 860
rect 499 820 504 825
rect 475 794 480 799
rect 479 783 484 788
rect 636 790 641 795
rect 607 589 612 594
rect 563 578 568 583
rect 629 573 634 578
rect 499 562 504 567
rect 479 510 484 515
rect 629 503 634 508
rect 605 481 610 486
<< metal2 >>
rect 477 1531 526 1534
rect 477 799 480 1064
rect 489 851 492 1100
rect 496 1079 499 1359
rect 503 1131 506 1384
rect 519 1172 522 1436
rect 558 1145 561 1482
rect 622 1406 647 1409
rect 575 1365 578 1383
rect 570 1362 578 1365
rect 612 1178 615 1389
rect 622 1366 625 1406
rect 601 1175 615 1178
rect 558 1142 571 1145
rect 519 892 522 1031
rect 601 1008 604 1175
rect 640 1075 643 1137
rect 563 1005 604 1008
rect 563 867 566 1005
rect 627 982 630 1064
rect 579 979 630 982
rect 481 515 484 783
rect 501 567 504 820
rect 520 747 523 751
rect 517 744 523 747
rect 517 608 520 744
rect 579 619 582 979
rect 636 795 639 855
rect 563 616 582 619
rect 563 583 566 616
rect 609 594 612 765
rect 607 486 610 589
rect 629 508 632 573
<< m123contact >>
rect 82 1666 87 1671
rect 523 1666 528 1671
rect 743 1664 748 1669
rect -15 1657 -10 1662
rect 2 1603 7 1608
rect 737 1586 742 1591
rect 599 1555 604 1560
rect -3 1395 2 1400
rect -3 1111 2 1116
rect -3 831 2 836
rect 522 1433 527 1438
rect 617 1419 622 1424
rect 599 1359 604 1364
rect 762 1392 767 1397
rect 546 1123 551 1128
rect 613 1153 618 1158
rect 611 1043 616 1048
rect 835 1013 840 1018
rect -22 548 -17 553
rect -3 547 2 552
rect 609 873 614 878
rect 609 765 614 770
rect 832 733 837 738
rect 559 559 564 564
rect 643 582 648 587
rect 713 583 718 588
rect 773 578 778 583
rect 643 573 648 578
rect 787 561 792 566
rect 700 482 705 487
rect 58 387 63 392
rect 809 387 814 392
<< metal3 >>
rect -13 1608 -10 1657
rect 83 1644 86 1666
rect -13 1605 2 1608
rect -13 1399 -10 1605
rect 59 1455 62 1580
rect 130 1513 133 1522
rect 524 1438 527 1666
rect 745 1630 748 1664
rect 745 1627 828 1630
rect 825 1625 828 1627
rect 601 1461 604 1555
rect 737 1474 740 1586
rect 802 1496 805 1561
rect 872 1496 875 1503
rect 802 1493 833 1496
rect 737 1471 765 1474
rect 601 1458 737 1461
rect 622 1420 634 1423
rect -13 1396 -3 1399
rect -13 1115 -10 1396
rect 631 1362 634 1420
rect 631 1359 654 1362
rect 59 1171 62 1301
rect 130 1229 133 1243
rect 600 1197 603 1359
rect 600 1194 616 1197
rect 613 1158 616 1194
rect 734 1162 737 1458
rect 762 1397 765 1471
rect 762 1185 765 1392
rect 830 1372 833 1493
rect 854 1493 875 1496
rect 854 1431 857 1493
rect 829 1304 832 1367
rect 829 1301 872 1304
rect 762 1182 839 1185
rect 734 1159 809 1162
rect -13 1112 -3 1115
rect -13 835 -10 1112
rect 59 891 62 1017
rect 130 949 133 959
rect -13 832 -3 835
rect -13 551 -10 832
rect 59 607 62 737
rect 130 665 133 679
rect 548 625 551 1123
rect 613 1048 616 1153
rect 611 878 614 1043
rect 610 770 613 873
rect 806 636 809 1159
rect 836 1018 839 1182
rect 869 1053 872 1301
rect 901 1243 904 1309
rect 901 1240 974 1243
rect 971 1099 974 1240
rect 835 994 838 1013
rect 713 633 809 636
rect 832 991 838 994
rect 832 738 835 991
rect 867 775 870 1029
rect 924 836 927 977
rect 924 833 971 836
rect 968 819 971 833
rect 866 773 870 775
rect 867 772 870 773
rect 845 751 864 754
rect 548 622 646 625
rect 643 587 646 622
rect 713 588 716 633
rect 832 620 835 733
rect 787 617 835 620
rect 643 562 646 573
rect 564 559 646 562
rect -17 548 -3 551
rect 778 542 781 581
rect 787 566 790 617
rect 702 539 781 542
rect 845 541 848 751
rect 921 681 924 697
rect 869 678 924 681
rect 869 600 872 678
rect 702 487 705 539
rect 810 524 815 529
rect 59 392 62 453
rect 810 392 813 524
use ffi  ffi_0
timestamp 1618618094
transform 1 0 16 0 -1 1613
box -14 -42 207 91
use ffipg  ffipg_0
timestamp 1618623899
transform 1 0 2 0 1 1243
box -4 0 470 271
use sumffo  sumffo_0
timestamp 1618628987
transform 1 0 618 0 -1 1627
box -3 -9 349 129
use nor  nor_0
timestamp 1618580541
transform 1 0 519 0 1 1397
box 0 -30 34 39
use inv  inv_0
timestamp 1618579805
transform 1 0 553 0 1 1390
box 0 -15 24 33
use nand  nand_0
timestamp 1618580231
transform 1 0 577 0 1 1396
box 0 -35 34 27
use sumffo  sumffo_1
timestamp 1618628987
transform 1 0 645 0 -1 1433
box -3 -9 349 129
use ffipg  ffipg_1
timestamp 1618623899
transform 1 0 2 0 1 959
box -4 0 470 271
use nand  nand_1
timestamp 1618580231
transform 1 0 579 0 -1 1134
box 0 -35 34 27
use inv  inv_2
timestamp 1618579805
transform 1 0 613 0 -1 1141
box 0 -15 24 33
use cla  cla_0
timestamp 1618627066
transform 1 0 516 0 1 1077
box -9 -46 112 95
use nor  nor_1
timestamp 1618580541
transform 1 0 648 0 1 1075
box 0 -30 34 39
use inv  inv_1
timestamp 1618579805
transform 1 0 682 0 1 1068
box 0 -15 24 33
use sumffo  sumffo_2
timestamp 1618628987
transform 1 0 717 0 1 975
box -3 -9 349 129
use ffipg  ffipg_2
timestamp 1618623899
transform 1 0 2 0 1 679
box -4 0 470 271
use nand  nand_2
timestamp 1618580231
transform 1 0 575 0 -1 854
box 0 -35 34 27
use inv  inv_3
timestamp 1618579805
transform 1 0 609 0 -1 861
box 0 -15 24 33
use cla  cla_1
timestamp 1618627066
transform 1 0 516 0 1 797
box -9 -46 112 95
use nor  nor_2
timestamp 1618580541
transform 1 0 647 0 1 795
box 0 -30 34 39
use inv  inv_4
timestamp 1618579805
transform 1 0 681 0 1 788
box 0 -15 24 33
use sumffo  sumffo_3
timestamp 1618628987
transform 1 0 714 0 1 695
box -3 -9 349 129
use ffipg  ffipg_3
timestamp 1618623899
transform 1 0 2 0 1 395
box -4 0 470 271
use nand  nand_3
timestamp 1618580231
transform 1 0 573 0 -1 570
box 0 -35 34 27
use inv  inv_5
timestamp 1618579805
transform 1 0 607 0 -1 577
box 0 -15 24 33
use nand  nand_4
timestamp 1618580231
transform 1 0 651 0 -1 574
box 0 -35 34 27
use inv  inv_7
timestamp 1618579805
transform 1 0 685 0 -1 581
box 0 -15 24 33
use nand  nand_5
timestamp 1618580231
transform 1 0 718 0 -1 575
box 0 -35 34 27
use inv  inv_8
timestamp 1618579805
transform 1 0 752 0 -1 582
box 0 -15 24 33
use cla  cla_2
timestamp 1618627066
transform 1 0 513 0 1 513
box -9 -46 112 95
use nor  nor_3
timestamp 1618580541
transform 1 0 638 0 1 508
box 0 -30 34 39
use inv  inv_6
timestamp 1618579805
transform 1 0 672 0 1 501
box 0 -15 24 33
use nor  nor_4
timestamp 1618580541
transform 1 0 705 0 1 495
box 0 -30 34 39
use inv  inv_9
timestamp 1618579805
transform 1 0 739 0 1 488
box 0 -15 24 33
use ffo  ffo_0
timestamp 1618618535
transform 1 0 801 0 -1 569
box -14 -42 207 91
<< labels >>
rlabel metal1 -17 1659 -17 1662 3 clk
rlabel metal1 -17 1666 -17 1669 4 vdd!
rlabel metal1 -2 387 -2 390 1 gnd!
rlabel metal1 -17 1552 -17 1555 3 cinin
rlabel metal1 -17 1273 -17 1276 3 y1in
rlabel metal1 -17 1480 -17 1483 3 x1in
rlabel metal1 -17 1196 -17 1199 3 x2in
rlabel metal1 -17 989 -17 992 3 y2in
rlabel metal1 -17 916 -17 919 3 x3in
rlabel metal1 -17 709 -17 712 3 y3in
rlabel metal1 -17 632 -17 635 3 x4in
rlabel metal1 -17 425 -17 428 3 y4in
rlabel metal1 1065 727 1065 730 7 z4o
rlabel metal1 1010 567 1010 570 1 couto
rlabel metal1 1068 1007 1068 1010 7 z3o
rlabel metal1 996 1398 996 1401 1 z2o
rlabel metal1 969 1592 969 1595 1 z1o
rlabel metal1 -24 548 -24 551 3 test
<< end >>
