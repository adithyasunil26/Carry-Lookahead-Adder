magic
tech scmos
timestamp 1618621484
<< metal1 >>
rect 3 109 118 111
rect 3 108 172 109
rect 3 74 6 108
rect 115 106 172 108
rect -1 70 0 73
rect 3 69 8 74
rect 115 59 118 106
rect 115 56 125 59
rect 119 50 125 53
rect -1 16 0 19
rect 3 15 8 20
rect 5 -3 8 15
rect 119 2 122 50
rect 169 39 172 106
rect 217 88 219 91
rect 217 61 219 64
rect 169 36 175 39
rect 209 35 219 38
rect 159 31 162 34
rect 141 25 144 31
rect 165 30 175 33
rect 165 2 168 30
rect 44 -1 168 2
rect 44 -3 47 -1
rect 5 -6 47 -3
<< m2contact >>
rect 156 53 161 58
rect 111 35 116 40
rect 212 86 217 91
rect 212 59 217 64
<< metal2 >>
rect 113 88 212 91
rect 3 69 8 74
rect 113 40 116 88
rect 165 61 212 64
rect 165 58 168 61
rect 161 55 168 58
rect 3 15 8 20
<< m123contact >>
rect 99 96 104 101
rect 139 97 144 102
rect 184 68 189 73
rect 140 20 145 25
rect 104 6 109 11
rect 177 6 182 11
<< metal3 >>
rect 104 98 139 101
rect 144 97 165 100
rect 162 71 165 97
rect 162 68 184 71
rect 141 9 144 20
rect 109 6 177 9
use xor  xor_0
timestamp 1618605809
transform 1 0 53 0 1 56
box -53 -56 59 49
use nor  nor_0
timestamp 1618580541
transform 1 0 125 0 1 61
box 0 -30 34 39
use nand  nand_0
timestamp 1618580231
transform 1 0 175 0 1 41
box 0 -35 34 27
<< labels >>
rlabel metal1 219 35 219 38 7 g
rlabel metal1 219 61 219 64 7 p
rlabel metal1 219 88 219 91 7 k
rlabel metal1 -1 70 -1 73 3 x
rlabel metal1 -1 16 -1 19 3 y
<< end >>
