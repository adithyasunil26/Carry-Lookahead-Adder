* SPICE3 file created from adder.ext - technology: scmos

.option scale=0.09u

M1000 nand_1/a_13_n26# cla_0/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=3510 ps=2284
M1001 vdd cin inv_2/in inv_2/w_0_6# pfet w=12 l=2
+  ad=7020 pd=3668 as=96 ps=40
M1002 inv_2/in cla_0/l vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 inv_2/in cin nand_1/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1004 nand_0/a_13_n26# inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1005 vdd cla_0/g0 nand_2/b nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1006 nand_2/b inv_0/op vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 nand_2/b cla_0/g0 nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1008 nand_2/a_13_n26# cla_1/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 vdd nand_2/b inv_3/in inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1010 inv_3/in cla_1/l vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 inv_3/in nand_2/b nand_2/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1012 nand_3/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1013 vdd cla_0/n inv_5/in inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1014 inv_5/in cla_2/l vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 inv_5/in cla_0/n nand_3/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1016 nand_4/a_13_n26# cla_2/l gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1017 vdd cla_0/l inv_7/in inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1018 inv_7/in cla_2/l vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 inv_7/in cla_0/l nand_4/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1020 cla_0/nand_0/a_13_n26# cla_0/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1021 vdd cla_1/g0 cla_0/n cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1022 cla_0/n cla_0/inv_0/op vdd cla_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 cla_0/n cla_1/g0 cla_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1024 cla_0/inv_0/op cla_0/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1025 cla_0/inv_0/op cla_0/inv_0/in vdd cla_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1026 cla_0/l nor_0/a cla_0/nor_0/a_13_6# cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1027 cla_0/nor_0/a_13_6# cla_1/p0 vdd cla_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 gnd nor_0/a cla_0/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1029 cla_0/l cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 cla_0/inv_0/in cla_0/g0 cla_0/nor_1/a_13_6# cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1031 cla_0/nor_1/a_13_6# cla_1/p0 vdd cla_0/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 gnd cla_0/g0 cla_0/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1033 cla_0/inv_0/in cla_1/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 nand_5/a_13_n26# inv_7/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1035 vdd cin inv_8/in inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1036 inv_8/in inv_7/op vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 inv_8/in cin nand_5/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1038 cla_1/nand_0/a_13_n26# cla_1/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1039 vdd cla_2/g0 cla_1/n cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1040 cla_1/n cla_1/inv_0/op vdd cla_1/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 cla_1/n cla_2/g0 cla_1/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1042 cla_1/inv_0/op cla_1/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1043 cla_1/inv_0/op cla_1/inv_0/in vdd cla_1/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1044 cla_1/l cla_1/p0 cla_1/nor_0/a_13_6# cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1045 cla_1/nor_0/a_13_6# cla_2/p0 vdd cla_1/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd cla_1/p0 cla_1/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1047 cla_1/l cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 cla_1/inv_0/in cla_1/g0 cla_1/nor_1/a_13_6# cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1049 cla_1/nor_1/a_13_6# cla_2/p0 vdd cla_1/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd cla_1/g0 cla_1/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1051 cla_1/inv_0/in cla_2/p0 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 cla_2/nand_0/a_13_n26# cla_2/inv_0/op gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1053 vdd cla_2/g1 cla_2/n cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1054 cla_2/n cla_2/inv_0/op vdd cla_2/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 cla_2/n cla_2/g1 cla_2/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1056 cla_2/inv_0/op cla_2/inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 cla_2/inv_0/op cla_2/inv_0/in vdd cla_2/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1058 cla_2/l cla_2/p0 cla_2/nor_0/a_13_6# cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1059 cla_2/nor_0/a_13_6# cla_2/p1 vdd cla_2/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 gnd cla_2/p0 cla_2/l Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1061 cla_2/l cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 cla_2/inv_0/in cla_2/g0 cla_2/nor_1/a_13_6# cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1063 cla_2/nor_1/a_13_6# cla_2/p1 vdd cla_2/nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 gnd cla_2/g0 cla_2/inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1065 cla_2/inv_0/in cla_2/p1 gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 sumffo_0/xor_0/inv_0/op ffipg_0/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1067 sumffo_0/xor_0/inv_0/op ffipg_0/k vdd sumffo_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1068 sumffo_0/xor_0/inv_1/op cin gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1069 sumffo_0/xor_0/inv_1/op cin vdd sumffo_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1070 vdd cin sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1071 s1 cin sumffo_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1072 gnd sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1073 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/inv_1/op s1 sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1074 sumffo_0/xor_0/a_10_n43# ffipg_0/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 sumffo_0/xor_0/a_38_n43# sumffo_0/xor_0/inv_0/op s1 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 sumffo_0/xor_0/a_10_10# ffipg_0/k vdd sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 s1 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 sumffo_2/xor_0/inv_0/op inv_1/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 sumffo_2/xor_0/inv_0/op inv_1/op vdd sumffo_2/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1080 sumffo_2/xor_0/inv_1/op sumffo_2/c gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1081 sumffo_2/xor_0/inv_1/op sumffo_2/c vdd sumffo_2/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1082 vdd sumffo_2/c sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1083 s3 sumffo_2/c sumffo_2/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1084 gnd sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1085 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/inv_1/op s3 sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1086 sumffo_2/xor_0/a_10_n43# inv_1/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 sumffo_2/xor_0/a_38_n43# sumffo_2/xor_0/inv_0/op s3 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 sumffo_2/xor_0/a_10_10# inv_1/op vdd sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 s3 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 sumffo_1/xor_0/inv_0/op ffipg_1/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1091 sumffo_1/xor_0/inv_0/op ffipg_1/k vdd sumffo_1/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1092 sumffo_1/xor_0/inv_1/op nand_2/b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1093 sumffo_1/xor_0/inv_1/op nand_2/b vdd sumffo_1/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1094 vdd nand_2/b sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1095 s2 nand_2/b sumffo_1/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1096 gnd sumffo_1/xor_0/inv_1/op sumffo_1/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1097 sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/inv_1/op s2 sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1098 sumffo_1/xor_0/a_10_n43# ffipg_1/k gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 sumffo_1/xor_0/a_38_n43# sumffo_1/xor_0/inv_0/op s2 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 sumffo_1/xor_0/a_10_10# ffipg_1/k vdd sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 s2 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/a_10_10# sumffo_1/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 sumffo_3/xor_0/inv_0/op inv_4/op gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1103 sumffo_3/xor_0/inv_0/op inv_4/op vdd sumffo_3/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1104 sumffo_3/xor_0/inv_1/op ffipg_3/k gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1105 sumffo_3/xor_0/inv_1/op ffipg_3/k vdd sumffo_3/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1106 vdd ffipg_3/k sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1107 s4 ffipg_3/k sumffo_3/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1108 gnd sumffo_3/xor_0/inv_1/op sumffo_3/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1109 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/inv_1/op s4 sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1110 sumffo_3/xor_0/a_10_n43# inv_4/op gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 sumffo_3/xor_0/a_38_n43# sumffo_3/xor_0/inv_0/op s4 Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 sumffo_3/xor_0/a_10_10# inv_4/op vdd sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 s4 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 inv_0/op inv_0/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 inv_0/op inv_0/in vdd nor_0/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1116 inv_1/op inv_1/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1117 inv_1/op inv_1/in vdd nor_1/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1118 nor_1/b inv_2/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1119 nor_1/b inv_2/in vdd inv_2/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1120 inv_0/in cinbar nor_0/a_13_6# nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1121 nor_0/a_13_6# nor_0/a vdd nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd cinbar inv_0/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1123 inv_0/in nor_0/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 nor_2/b inv_3/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1125 nor_2/b inv_3/in vdd inv_3/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1126 inv_1/in nor_1/b nor_1/a_13_6# nor_1/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1127 nor_1/a_13_6# cla_0/n vdd nor_1/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 gnd nor_1/b inv_1/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1129 inv_1/in cla_0/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 inv_4/op inv_4/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1131 inv_4/op inv_4/in vdd nor_2/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1132 inv_4/in nor_2/b nor_2/a_13_6# nor_2/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1133 nor_2/a_13_6# cla_1/n vdd nor_2/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd nor_2/b inv_4/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1135 inv_4/in cla_1/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 nor_4/b inv_6/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1137 nor_4/b inv_6/in vdd nor_3/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1138 inv_6/in nor_3/b nor_3/a_13_6# nor_3/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1139 nor_3/a_13_6# cla_2/n vdd nor_3/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd nor_3/b inv_6/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1141 inv_6/in cla_2/n gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 nor_3/b inv_5/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1143 nor_3/b inv_5/in vdd inv_5/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1144 inv_9/in nor_4/b nor_4/a_13_6# nor_4/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1145 nor_4/a_13_6# nor_4/a vdd nor_4/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 gnd nor_4/b inv_9/in Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1147 inv_9/in nor_4/a gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 inv_7/op inv_7/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1149 inv_7/op inv_7/in vdd inv_7/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1150 nor_4/a inv_8/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1151 nor_4/a inv_8/in vdd inv_8/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1152 ffipg_0/pggen_0/nand_0/a_13_n26# x1in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1153 vdd y1in cla_0/g0 ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1154 cla_0/g0 x1in vdd ffipg_0/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 cla_0/g0 y1in ffipg_0/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1156 ffipg_0/pggen_0/xor_0/inv_0/op x1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1157 ffipg_0/pggen_0/xor_0/inv_0/op x1in vdd ffipg_0/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1158 ffipg_0/pggen_0/xor_0/inv_1/op y1in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1159 ffipg_0/pggen_0/xor_0/inv_1/op y1in vdd ffipg_0/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1160 vdd y1in ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1161 ffipg_0/k y1in ffipg_0/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1162 gnd ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1163 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/inv_1/op ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1164 ffipg_0/pggen_0/xor_0/a_10_n43# x1in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ffipg_0/pggen_0/xor_0/a_38_n43# ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 ffipg_0/pggen_0/xor_0/a_10_10# x1in vdd ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 nor_0/a x1in ffipg_0/pggen_0/nor_0/a_13_6# ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1169 ffipg_0/pggen_0/nor_0/a_13_6# y1in vdd ffipg_0/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 gnd x1in nor_0/a Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1171 nor_0/a y1in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 cout inv_9/in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1173 cout inv_9/in vdd nor_4/w_0_0# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1174 ffipg_1/pggen_0/nand_0/a_13_n26# x2in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1175 vdd y2in cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1176 cla_1/g0 x2in vdd ffipg_1/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 cla_1/g0 y2in ffipg_1/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1178 ffipg_1/pggen_0/xor_0/inv_0/op x2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1179 ffipg_1/pggen_0/xor_0/inv_0/op x2in vdd ffipg_1/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1180 ffipg_1/pggen_0/xor_0/inv_1/op y2in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1181 ffipg_1/pggen_0/xor_0/inv_1/op y2in vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1182 vdd y2in ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1183 ffipg_1/k y2in ffipg_1/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1184 gnd ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1185 ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1186 ffipg_1/pggen_0/xor_0/a_10_n43# x2in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 ffipg_1/pggen_0/xor_0/a_38_n43# ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ffipg_1/pggen_0/xor_0/a_10_10# x2in vdd ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op ffipg_1/pggen_0/xor_0/a_10_10# ffipg_1/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 cla_1/p0 x2in ffipg_1/pggen_0/nor_0/a_13_6# ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1191 ffipg_1/pggen_0/nor_0/a_13_6# y2in vdd ffipg_1/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 gnd x2in cla_1/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1193 cla_1/p0 y2in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ffipg_2/pggen_0/nand_0/a_13_n26# x3in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1195 vdd y3in cla_2/g0 ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1196 cla_2/g0 x3in vdd ffipg_2/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 cla_2/g0 y3in ffipg_2/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1198 ffipg_2/pggen_0/xor_0/inv_0/op x3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1199 ffipg_2/pggen_0/xor_0/inv_0/op x3in vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1200 ffipg_2/pggen_0/xor_0/inv_1/op y3in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1201 ffipg_2/pggen_0/xor_0/inv_1/op y3in vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1202 vdd y3in ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1203 ffipg_2/k y3in ffipg_2/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1204 gnd ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1205 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1206 ffipg_2/pggen_0/xor_0/a_10_n43# x3in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ffipg_2/pggen_0/xor_0/a_38_n43# ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 ffipg_2/pggen_0/xor_0/a_10_10# x3in vdd ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 ffipg_2/k ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 cla_2/p0 x3in ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1211 ffipg_2/pggen_0/nor_0/a_13_6# y3in vdd ffipg_2/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 gnd x3in cla_2/p0 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1213 cla_2/p0 y3in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 ffipg_3/pggen_0/nand_0/a_13_n26# x4in gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1215 vdd y4in cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1216 cla_2/g1 x4in vdd ffipg_3/pggen_0/nand_0/w_0_0# pfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 cla_2/g1 y4in ffipg_3/pggen_0/nand_0/a_13_n26# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1218 ffipg_3/pggen_0/xor_0/inv_0/op x4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1219 ffipg_3/pggen_0/xor_0/inv_0/op x4in vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1220 ffipg_3/pggen_0/xor_0/inv_1/op y4in gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1221 ffipg_3/pggen_0/xor_0/inv_1/op y4in vdd ffipg_3/pggen_0/xor_0/inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1222 vdd y4in ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=432 ps=180
M1223 ffipg_3/k y4in ffipg_3/pggen_0/xor_0/a_10_n43# Gnd nfet w=12 l=2
+  ad=120 pd=68 as=96 ps=40
M1224 gnd ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/pggen_0/xor_0/a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1225 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/inv_1/op ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=192 ps=64
M1226 ffipg_3/pggen_0/xor_0/a_10_n43# x4in gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ffipg_3/pggen_0/xor_0/a_38_n43# ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/k Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ffipg_3/pggen_0/xor_0/a_10_10# x4in vdd ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 cla_2/p1 x4in ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=120 pd=58 as=192 ps=64
M1231 ffipg_3/pggen_0/nor_0/a_13_6# y4in vdd ffipg_3/pggen_0/nor_0/w_0_0# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 gnd x4in cla_2/p1 Gnd nfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1233 cla_2/p1 y4in gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 ffipg_2/pggen_0/nand_0/w_0_0# x3in 0.06fF
C1 gnd cla_1/nand_0/a_13_n26# 0.01fF
C2 cout vdd 0.15fF
C3 gnd s1 0.14fF
C4 s3 cin 0.28fF
C5 ffipg_1/pggen_0/xor_0/a_10_10# vdd 0.93fF
C6 inv_4/op inv_4/in 0.04fF
C7 sumffo_1/xor_0/inv_1/op s2 0.52fF
C8 nor_0/w_0_0# vdd 0.46fF
C9 ffipg_1/pggen_0/xor_0/inv_0/op x2in 0.27fF
C10 y2in cla_1/p0 0.03fF
C11 nor_0/w_0_0# cin 0.16fF
C12 ffipg_0/k ffipg_0/pggen_0/xor_0/a_10_10# 0.45fF
C13 cla_1/g0 ffipg_1/pggen_0/nand_0/w_0_0# 0.04fF
C14 ffipg_3/k vdd 0.35fF
C15 cla_1/g0 cla_0/n 0.13fF
C16 gnd ffipg_0/pggen_0/xor_0/inv_1/op 0.20fF
C17 vdd ffipg_1/pggen_0/nand_0/w_0_0# 0.10fF
C18 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/a_10_10# 0.16fF
C19 cla_2/g0 cla_1/nand_0/w_0_0# 0.06fF
C20 ffipg_0/k cinbar 0.06fF
C21 gnd cla_1/l 0.18fF
C22 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/inv_0/w_0_6# 0.03fF
C23 cla_0/n vdd 0.56fF
C24 sumffo_1/xor_0/inv_0/op sumffo_1/xor_0/inv_1/op 0.08fF
C25 ffipg_0/pggen_0/xor_0/inv_0/op vdd 0.15fF
C26 gnd cla_2/inv_0/in 0.30fF
C27 gnd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.02fF
C28 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_1/op 0.52fF
C29 inv_3/in inv_3/w_0_6# 0.10fF
C30 cla_2/p1 vdd 0.31fF
C31 nor_4/b nor_4/w_0_0# 0.06fF
C32 cla_2/g0 y3in 0.13fF
C33 sumffo_1/xor_0/w_n3_4# nand_2/b 0.06fF
C34 cout inv_9/in 0.04fF
C35 y2in ffipg_1/pggen_0/xor_0/a_10_10# 0.12fF
C36 cla_0/n inv_5/w_0_6# 0.06fF
C37 nor_0/a y1in 0.03fF
C38 gnd ffipg_2/k 0.14fF
C39 cla_1/g0 nand_2/b 0.06fF
C40 ffipg_0/pggen_0/nor_0/w_0_0# ffipg_0/k 0.21fF
C41 inv_1/op sumffo_2/c 0.09fF
C42 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/xor_0/inv_1/op 0.03fF
C43 ffipg_1/pggen_0/xor_0/inv_1/op x2in 0.06fF
C44 cla_2/g0 cla_2/p0 0.08fF
C45 nand_2/b vdd 0.92fF
C46 cin sumffo_2/xor_0/a_38_n43# 0.01fF
C47 cla_0/l inv_3/w_0_6# 0.00fF
C48 gnd inv_3/in 0.17fF
C49 nand_2/b cin 0.04fF
C50 cla_0/inv_0/w_0_6# vdd 0.06fF
C51 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C52 y2in ffipg_1/pggen_0/nand_0/w_0_0# 0.06fF
C53 vdd y4in 0.10fF
C54 nor_3/w_0_0# vdd 0.14fF
C55 sumffo_1/xor_0/inv_0/w_0_6# ffipg_1/k 0.06fF
C56 inv_2/w_0_6# nor_1/b 0.03fF
C57 sumffo_2/xor_0/inv_0/w_0_6# sumffo_2/xor_0/inv_0/op 0.03fF
C58 gnd x3in 0.31fF
C59 gnd cla_2/l 0.24fF
C60 cla_2/g0 ffipg_3/k 0.06fF
C61 gnd cla_0/g0 0.70fF
C62 cla_1/inv_0/op vdd 0.17fF
C63 cla_0/l inv_7/in 0.13fF
C64 cla_1/g0 cla_1/nor_1/w_0_0# 0.06fF
C65 cla_2/g0 cla_0/n 0.06fF
C66 inv_4/op sumffo_3/xor_0/w_n3_4# 0.06fF
C67 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# x1in 0.06fF
C68 gnd x2in 0.31fF
C69 gnd cla_0/l 0.98fF
C70 cla_2/g0 cla_2/p1 0.30fF
C71 cla_1/nor_1/w_0_0# vdd 0.31fF
C72 cla_2/g1 cla_2/nor_1/w_0_0# 0.02fF
C73 gnd ffipg_2/pggen_0/xor_0/w_n3_4# 0.02fF
C74 gnd sumffo_0/xor_0/inv_1/op 0.20fF
C75 nor_0/a vdd 0.35fF
C76 cla_0/n inv_5/in 0.13fF
C77 ffipg_0/pggen_0/xor_0/a_10_10# y1in 0.12fF
C78 sumffo_1/xor_0/inv_0/op s2 0.06fF
C79 ffipg_0/k sumffo_0/xor_0/inv_1/op 0.06fF
C80 cla_2/nor_0/w_0_0# vdd 0.31fF
C81 cla_1/g0 cla_0/inv_0/in 0.04fF
C82 x4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C83 sumffo_1/xor_0/inv_1/w_0_6# sumffo_1/xor_0/inv_1/op 0.03fF
C84 cla_0/inv_0/in vdd 0.05fF
C85 ffipg_1/k cla_0/g0 0.06fF
C86 gnd cla_0/inv_0/op 0.10fF
C87 cla_1/p0 cla_0/nor_1/w_0_0# 0.06fF
C88 nor_0/w_0_0# inv_0/op 0.10fF
C89 y1in ffipg_0/pggen_0/xor_0/inv_1/op 0.22fF
C90 inv_4/op nor_2/w_0_0# 0.03fF
C91 ffipg_1/k x2in 0.46fF
C92 cla_2/inv_0/w_0_6# vdd 0.06fF
C93 nor_1/w_0_0# vdd 0.17fF
C94 gnd ffipg_2/pggen_0/xor_0/inv_0/op 0.21fF
C95 inv_4/op gnd 0.32fF
C96 y3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C97 inv_1/in cla_0/n 0.02fF
C98 gnd sumffo_1/xor_0/inv_1/op 0.20fF
C99 nor_4/b vdd 0.15fF
C100 cla_0/l cla_0/nor_0/w_0_0# 0.05fF
C101 ffipg_3/pggen_0/xor_0/inv_0/op vdd 0.15fF
C102 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C103 sumffo_1/xor_0/a_10_10# s2 0.45fF
C104 cla_1/inv_0/w_0_6# vdd 0.06fF
C105 y3in ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C106 cla_2/p0 cla_1/p0 0.24fF
C107 ffipg_0/pggen_0/nor_0/w_0_0# y1in 0.06fF
C108 sumffo_2/xor_0/inv_0/w_0_6# vdd 0.09fF
C109 cla_2/g0 cla_1/inv_0/op 0.35fF
C110 cla_2/p0 y3in 0.03fF
C111 gnd inv_2/w_0_6# 0.02fF
C112 nor_2/b inv_3/in 0.04fF
C113 s3 sumffo_2/xor_0/inv_1/op 0.52fF
C114 cla_2/p0 ffipg_2/pggen_0/nor_0/w_0_0# 0.05fF
C115 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C116 gnd sumffo_2/c 0.15fF
C117 gnd cla_0/nand_0/w_0_0# 0.01fF
C118 cla_2/g0 cla_1/nor_1/w_0_0# 0.02fF
C119 ffipg_0/pggen_0/xor_0/a_10_10# vdd 0.93fF
C120 ffipg_3/k sumffo_3/xor_0/inv_1/op 0.22fF
C121 ffipg_3/k ffipg_3/pggen_0/xor_0/w_n3_4# 0.02fF
C122 inv_4/in cla_1/n 0.02fF
C123 gnd inv_0/in 0.24fF
C124 sumffo_2/xor_0/a_10_10# sumffo_2/xor_0/w_n3_4# 0.16fF
C125 sumffo_0/xor_0/inv_1/w_0_6# vdd 0.07fF
C126 ffipg_1/k sumffo_1/xor_0/inv_1/op 0.06fF
C127 cla_2/l inv_7/w_0_6# 0.06fF
C128 x4in ffipg_3/k 0.46fF
C129 nor_3/w_0_0# nor_3/b 0.06fF
C130 cinbar vdd 0.16fF
C131 sumffo_0/xor_0/inv_1/w_0_6# cin 0.23fF
C132 cla_1/p0 ffipg_1/pggen_0/nand_0/w_0_0# 0.24fF
C133 ffipg_3/pggen_0/nor_0/w_0_0# vdd 0.11fF
C134 vdd ffipg_0/pggen_0/xor_0/inv_1/op 0.15fF
C135 sumffo_3/xor_0/a_38_n43# cin 0.01fF
C136 nor_4/b inv_9/in 0.16fF
C137 cla_1/l vdd 0.22fF
C138 cla_0/l inv_7/w_0_6# 0.06fF
C139 x4in cla_2/p1 0.22fF
C140 inv_2/in inv_2/w_0_6# 0.10fF
C141 cla_0/g0 y1in 0.13fF
C142 cla_2/inv_0/in vdd 0.05fF
C143 vdd ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C144 inv_6/in cla_2/n 0.02fF
C145 ffipg_1/k ffipg_1/pggen_0/nor_0/w_0_0# 0.21fF
C146 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/k 0.52fF
C147 sumffo_1/xor_0/inv_0/w_0_6# vdd 0.09fF
C148 s4 sumffo_3/xor_0/w_n3_4# 0.02fF
C149 ffipg_0/pggen_0/nand_0/w_0_0# nor_0/a 0.24fF
C150 gnd x1in 0.22fF
C151 cla_2/p0 ffipg_3/k 0.06fF
C152 ffipg_0/pggen_0/nor_0/w_0_0# vdd 0.11fF
C153 cla_1/g0 ffipg_2/k 0.06fF
C154 cla_2/g1 ffipg_3/pggen_0/nand_0/w_0_0# 0.04fF
C155 ffipg_0/k x1in 0.46fF
C156 vdd ffipg_2/k 0.25fF
C157 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# ffipg_3/pggen_0/xor_0/inv_1/op 0.03fF
C158 gnd inv_6/in 0.24fF
C159 cla_2/p0 cla_2/p1 0.24fF
C160 y4in ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C161 inv_3/in vdd 0.30fF
C162 gnd s2 0.14fF
C163 vdd ffipg_3/pggen_0/xor_0/a_10_10# 0.93fF
C164 inv_4/in nor_2/w_0_0# 0.11fF
C165 x4in y4in 0.73fF
C166 ffipg_2/pggen_0/xor_0/inv_1/op x3in 0.06fF
C167 gnd inv_4/in 0.24fF
C168 ffipg_1/pggen_0/xor_0/inv_1/op ffipg_1/pggen_0/xor_0/inv_0/op 0.08fF
C169 sumffo_2/xor_0/a_10_10# vdd 0.93fF
C170 gnd s4 0.14fF
C171 cla_1/nand_0/w_0_0# cla_1/inv_0/op 0.06fF
C172 cla_0/n ffipg_3/k 0.06fF
C173 inv_4/op sumffo_3/xor_0/inv_0/op 0.27fF
C174 cla_1/g0 cla_0/g0 0.14fF
C175 sumffo_3/xor_0/inv_1/w_0_6# vdd 0.06fF
C176 vdd x3in 0.93fF
C177 inv_1/in nor_1/w_0_0# 0.11fF
C178 ffipg_3/k cla_2/p1 0.05fF
C179 cin sumffo_2/xor_0/a_10_10# 0.04fF
C180 sumffo_0/xor_0/w_n3_4# s1 0.02fF
C181 cla_2/l vdd 0.38fF
C182 sumffo_2/c sumffo_2/xor_0/inv_0/op 0.20fF
C183 cla_0/g0 vdd 0.53fF
C184 gnd sumffo_1/xor_0/inv_0/op 0.17fF
C185 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C186 cla_0/l cla_1/g0 0.12fF
C187 cin cla_0/g0 0.08fF
C188 cla_2/g1 cla_2/nand_0/w_0_0# 0.06fF
C189 sumffo_2/c sumffo_2/xor_0/w_n3_4# 0.06fF
C190 cla_2/inv_0/w_0_6# cla_2/inv_0/op 0.03fF
C191 vdd x2in 0.93fF
C192 cla_2/g0 cla_2/inv_0/in 0.16fF
C193 nor_0/w_0_0# nand_2/b 0.04fF
C194 gnd inv_1/op 0.32fF
C195 cla_0/l vdd 0.53fF
C196 sumffo_0/xor_0/inv_0/op s1 0.06fF
C197 cla_1/p0 nor_0/a 0.24fF
C198 cla_2/l inv_5/w_0_6# 0.08fF
C199 ffipg_2/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C200 sumffo_3/xor_0/a_10_10# s4 0.45fF
C201 gnd cla_1/inv_0/in 0.30fF
C202 cla_0/l cin 0.33fF
C203 sumffo_0/xor_0/inv_1/op vdd 0.15fF
C204 gnd ffipg_3/pggen_0/xor_0/inv_1/op 0.20fF
C205 sumffo_0/xor_0/inv_1/op cin 0.22fF
C206 gnd ffipg_1/pggen_0/xor_0/inv_0/op 0.21fF
C207 cla_0/inv_0/in cla_1/p0 0.02fF
C208 cla_1/g0 cla_0/inv_0/op 0.35fF
C209 cla_2/nand_0/w_0_0# cla_2/n 0.04fF
C210 cla_0/inv_0/in cla_0/nor_1/w_0_0# 0.05fF
C211 nand_2/b cla_0/n 0.06fF
C212 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_0/op 0.08fF
C213 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_1/op 0.06fF
C214 ffipg_3/k y4in 0.07fF
C215 ffipg_1/pggen_0/xor_0/w_n3_4# x2in 0.06fF
C216 cla_0/inv_0/op vdd 0.17fF
C217 ffipg_0/pggen_0/xor_0/a_10_10# ffipg_0/pggen_0/xor_0/w_n3_4# 0.16fF
C218 ffipg_1/k sumffo_1/xor_0/inv_0/op 0.27fF
C219 cla_2/p0 cla_1/nor_1/w_0_0# 0.06fF
C220 gnd nor_1/b 0.10fF
C221 ffipg_2/pggen_0/xor_0/inv_0/op vdd 0.15fF
C222 inv_4/op vdd 0.26fF
C223 cla_2/p1 y4in 0.03fF
C224 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/w_n3_4# 0.06fF
C225 cla_2/g1 cla_2/n 0.13fF
C226 cla_2/p0 cla_2/nor_0/w_0_0# 0.06fF
C227 nor_2/w_0_0# cla_1/n 0.06fF
C228 gnd cla_2/nand_0/w_0_0# 0.08fF
C229 ffipg_0/pggen_0/xor_0/w_n3_4# ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C230 y2in x2in 0.73fF
C231 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# y1in 0.23fF
C232 nor_0/w_0_0# nor_0/a 0.06fF
C233 sumffo_1/xor_0/inv_1/op vdd 0.15fF
C234 gnd cla_1/n 0.24fF
C235 x4in ffipg_3/pggen_0/xor_0/inv_0/op 0.27fF
C236 cla_0/n cla_1/inv_0/op 0.06fF
C237 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C238 cla_2/nor_1/w_0_0# vdd 0.31fF
C239 x1in y1in 0.73fF
C240 cin sumffo_1/xor_0/inv_1/op 0.04fF
C241 cla_1/nor_0/w_0_0# vdd 0.31fF
C242 cla_2/inv_0/in cla_2/inv_0/op 0.04fF
C243 cla_2/g1 gnd 0.30fF
C244 inv_2/w_0_6# vdd 0.15fF
C245 cla_0/nand_0/w_0_0# cla_1/g0 0.06fF
C246 inv_2/in nor_1/b 0.04fF
C247 sumffo_2/c vdd 0.10fF
C248 cla_2/g0 cla_0/l 0.05fF
C249 inv_4/in nor_2/b 0.16fF
C250 inv_2/w_0_6# cin 0.06fF
C251 cla_2/l inv_5/in 0.05fF
C252 gnd ffipg_1/pggen_0/xor_0/inv_1/op 0.24fF
C253 cla_0/nand_0/w_0_0# vdd 0.10fF
C254 vdd ffipg_1/pggen_0/nor_0/w_0_0# 0.11fF
C255 gnd inv_3/w_0_6# 0.02fF
C256 inv_0/in vdd 0.07fF
C257 nor_4/a gnd 0.21fF
C258 cla_2/nor_0/w_0_0# cla_2/p1 0.06fF
C259 inv_4/op sumffo_3/xor_0/inv_0/w_0_6# 0.06fF
C260 inv_0/in cin 0.07fF
C261 x4in ffipg_3/pggen_0/nor_0/w_0_0# 0.06fF
C262 gnd cla_2/n 0.32fF
C263 ffipg_0/pggen_0/nand_0/a_13_n26# vdd 0.01fF
C264 ffipg_0/pggen_0/nand_0/w_0_0# cla_0/g0 0.04fF
C265 cla_1/p0 cla_1/l 0.16fF
C266 sumffo_3/xor_0/inv_0/op s4 0.06fF
C267 inv_1/op sumffo_2/xor_0/inv_0/op 0.27fF
C268 sumffo_0/xor_0/a_10_10# vdd 0.93fF
C269 x3in ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C270 x4in ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.06fF
C271 cla_2/l nor_3/b 0.10fF
C272 cla_0/n nor_1/w_0_0# 0.06fF
C273 sumffo_3/xor_0/a_10_10# sumffo_3/xor_0/w_n3_4# 0.16fF
C274 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/w_n3_4# 0.06fF
C275 sumffo_0/xor_0/a_10_10# cin 0.12fF
C276 inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C277 gnd inv_7/in 0.13fF
C278 vdd ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C279 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_0/op 0.06fF
C280 ffipg_1/k ffipg_1/pggen_0/xor_0/inv_1/op 0.52fF
C281 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C282 vdd x1in 0.97fF
C283 sumffo_1/xor_0/w_n3_4# s2 0.02fF
C284 cin sumffo_1/xor_0/a_38_n43# 0.01fF
C285 cla_1/inv_0/w_0_6# cla_0/n 0.26fF
C286 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_0/op 0.08fF
C287 inv_0/op cla_0/g0 0.32fF
C288 vdd ffipg_2/pggen_0/nand_0/a_13_n26# 0.01fF
C289 ffipg_0/k gnd 0.41fF
C290 cla_1/p0 ffipg_2/k 0.06fF
C291 y2in ffipg_1/pggen_0/nor_0/w_0_0# 0.06fF
C292 cla_2/p0 cla_1/l 0.02fF
C293 cla_2/g0 cla_2/nor_1/w_0_0# 0.06fF
C294 ffipg_3/pggen_0/xor_0/a_10_10# ffipg_3/pggen_0/xor_0/w_n3_4# 0.16fF
C295 y3in ffipg_2/k 0.07fF
C296 nor_4/a inv_8/w_0_6# 0.03fF
C297 inv_6/in vdd 0.09fF
C298 nor_0/w_0_0# cinbar 0.06fF
C299 ffipg_2/k ffipg_2/pggen_0/nor_0/w_0_0# 0.21fF
C300 cla_0/inv_0/in cla_0/inv_0/w_0_6# 0.06fF
C301 nor_4/a nor_4/w_0_0# 0.07fF
C302 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/inv_0/op 0.06fF
C303 sumffo_3/xor_0/inv_1/w_0_6# sumffo_3/xor_0/inv_1/op 0.03fF
C304 inv_4/in vdd 0.09fF
C305 cin s2 0.27fF
C306 ffipg_3/k ffipg_3/pggen_0/nor_0/w_0_0# 0.21fF
C307 nor_2/b cla_1/n 0.39fF
C308 gnd ffipg_1/k 0.39fF
C309 inv_2/in gnd 0.17fF
C310 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C311 cla_2/p0 ffipg_2/k 0.05fF
C312 y2in ffipg_1/pggen_0/xor_0/inv_1/w_0_6# 0.23fF
C313 sumffo_2/xor_0/inv_1/w_0_6# sumffo_2/c 0.23fF
C314 cla_0/g0 cla_1/p0 0.38fF
C315 y3in x3in 0.73fF
C316 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_1/op 0.08fF
C317 cla_0/g0 cla_0/nor_1/w_0_0# 0.06fF
C318 cin s4 0.16fF
C319 cla_0/n cla_1/l 0.07fF
C320 ffipg_3/pggen_0/nor_0/w_0_0# cla_2/p1 0.05fF
C321 x3in ffipg_2/pggen_0/nor_0/w_0_0# 0.06fF
C322 ffipg_3/pggen_0/xor_0/inv_0/op y4in 0.20fF
C323 cla_0/l cla_1/nand_0/w_0_0# 0.01fF
C324 nor_4/b nor_3/w_0_0# 0.03fF
C325 nor_4/a inv_8/in 0.04fF
C326 sumffo_1/xor_0/inv_0/op vdd 0.15fF
C327 vdd ffipg_2/pggen_0/xor_0/a_10_10# 0.93fF
C328 cla_1/p0 x2in 0.22fF
C329 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C330 cla_2/inv_0/in cla_2/p1 0.02fF
C331 vdd ffipg_3/pggen_0/nand_0/w_0_0# 0.10fF
C332 cla_0/l cla_1/p0 0.02fF
C333 cin sumffo_1/xor_0/inv_0/op 0.06fF
C334 inv_1/op vdd 0.26fF
C335 cla_1/g0 cla_1/inv_0/in 0.16fF
C336 nor_2/b inv_3/w_0_6# 0.03fF
C337 sumffo_1/xor_0/w_n3_4# sumffo_1/xor_0/a_10_10# 0.16fF
C338 s3 sumffo_2/xor_0/a_10_10# 0.45fF
C339 cla_1/inv_0/w_0_6# cla_1/inv_0/op 0.03fF
C340 cla_1/inv_0/in vdd 0.05fF
C341 y3in ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C342 cla_2/p0 x3in 0.22fF
C343 vdd ffipg_3/pggen_0/xor_0/inv_1/op 0.15fF
C344 cla_2/p0 cla_2/l 0.16fF
C345 sumffo_0/xor_0/a_10_10# sumffo_0/xor_0/w_n3_4# 0.16fF
C346 ffipg_0/k ffipg_0/pggen_0/nor_0/a_13_6# 0.01fF
C347 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/w_n3_4# 0.06fF
C348 vdd ffipg_1/pggen_0/xor_0/inv_0/op 0.15fF
C349 ffipg_2/pggen_0/nand_0/w_0_0# vdd 0.10fF
C350 gnd inv_8/in 0.13fF
C351 ffipg_3/k ffipg_3/pggen_0/xor_0/a_10_10# 0.45fF
C352 nand_2/b cla_1/l 0.31fF
C353 inv_4/op sumffo_3/xor_0/inv_1/op 0.06fF
C354 sumffo_1/xor_0/a_10_10# vdd 0.93fF
C355 nor_0/w_0_0# cla_0/g0 0.06fF
C356 ffipg_3/pggen_0/nor_0/w_0_0# y4in 0.06fF
C357 inv_7/w_0_6# inv_7/in 0.10fF
C358 vdd nor_1/b 0.25fF
C359 gnd sumffo_2/xor_0/inv_0/op 0.17fF
C360 sumffo_1/xor_0/a_10_10# cin 0.06fF
C361 nor_2/w_0_0# nor_2/b 0.06fF
C362 inv_0/op inv_0/in 0.04fF
C363 ffipg_3/k sumffo_3/xor_0/inv_1/w_0_6# 0.23fF
C364 ffipg_2/pggen_0/xor_0/inv_0/op y3in 0.20fF
C365 gnd nor_2/b 0.10fF
C366 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_0/op 0.06fF
C367 cla_2/nand_0/w_0_0# vdd 0.10fF
C368 inv_7/in inv_7/op 0.04fF
C369 ffipg_1/pggen_0/nand_0/a_13_n26# vdd 0.01fF
C370 ffipg_0/pggen_0/nand_0/w_0_0# x1in 0.06fF
C371 vdd cla_1/n 0.28fF
C372 cla_0/n cla_2/l 0.32fF
C373 gnd y1in 1.62fF
C374 gnd inv_7/op 0.10fF
C375 cla_2/l cla_2/p1 0.02fF
C376 cla_1/p0 cla_1/nor_0/w_0_0# 0.06fF
C377 cla_0/l ffipg_3/k 0.04fF
C378 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# vdd 0.06fF
C379 gnd sumffo_3/xor_0/inv_0/op 0.17fF
C380 ffipg_1/pggen_0/nand_0/w_0_0# x2in 0.06fF
C381 ffipg_0/k y1in 0.07fF
C382 nand_2/b inv_3/in 0.13fF
C383 cla_0/l cla_0/n 0.05fF
C384 cinbar nor_0/a 0.32fF
C385 cla_2/g1 vdd 0.35fF
C386 inv_8/w_0_6# inv_8/in 0.10fF
C387 y2in ffipg_1/pggen_0/xor_0/inv_0/op 0.20fF
C388 x1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C389 nor_3/b inv_6/in 0.16fF
C390 cla_1/p0 ffipg_1/pggen_0/nor_0/w_0_0# 0.05fF
C391 sumffo_2/xor_0/inv_1/op sumffo_2/c 0.22fF
C392 vdd ffipg_1/pggen_0/xor_0/inv_1/op 0.15fF
C393 vdd sumffo_3/xor_0/w_n3_4# 0.12fF
C394 ffipg_3/pggen_0/xor_0/a_10_10# y4in 0.12fF
C395 inv_3/w_0_6# vdd 0.15fF
C396 cla_2/g0 cla_1/inv_0/in 0.04fF
C397 cin sumffo_3/xor_0/w_n3_4# 0.01fF
C398 nor_4/a vdd 0.19fF
C399 sumffo_1/xor_0/inv_1/w_0_6# vdd 0.06fF
C400 cla_2/p0 cla_1/nor_0/w_0_0# 0.06fF
C401 nand_2/b cla_0/g0 0.13fF
C402 vdd cla_2/n 0.28fF
C403 cla_2/g0 ffipg_2/pggen_0/nand_0/w_0_0# 0.04fF
C404 ffipg_0/pggen_0/nor_0/w_0_0# nor_0/a 0.05fF
C405 inv_4/op ffipg_3/k 0.09fF
C406 cla_0/l nand_2/b 0.08fF
C407 gnd ffipg_2/pggen_0/xor_0/inv_1/op 0.24fF
C408 ffipg_1/pggen_0/xor_0/w_n3_4# ffipg_1/pggen_0/xor_0/inv_1/op 0.06fF
C409 inv_8/w_0_6# inv_7/op 0.06fF
C410 cla_2/inv_0/w_0_6# cla_2/inv_0/in 0.06fF
C411 inv_7/in vdd 0.30fF
C412 cla_0/l cla_0/inv_0/w_0_6# 0.00fF
C413 gnd cla_1/g0 0.28fF
C414 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# x2in 0.06fF
C415 nor_2/w_0_0# vdd 0.17fF
C416 gnd vdd 3.73fF
C417 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C418 cla_2/g0 cla_1/n 0.13fF
C419 inv_1/op inv_1/in 0.04fF
C420 nor_0/w_0_0# inv_0/in 0.11fF
C421 cla_2/nor_1/w_0_0# cla_2/p1 0.06fF
C422 gnd cin 0.74fF
C423 y2in ffipg_1/pggen_0/xor_0/inv_1/op 0.22fF
C424 ffipg_0/k vdd 0.33fF
C425 nand_2/b cla_0/inv_0/op 0.09fF
C426 sumffo_1/xor_0/w_n3_4# ffipg_1/k 0.06fF
C427 cla_0/l cla_1/inv_0/op 0.05fF
C428 ffipg_0/k cin 0.19fF
C429 cla_0/n sumffo_2/c 0.06fF
C430 nor_4/a inv_9/in 0.02fF
C431 gnd inv_5/w_0_6# 0.26fF
C432 cla_0/inv_0/w_0_6# cla_0/inv_0/op 0.03fF
C433 cla_0/g0 nor_0/a 0.57fF
C434 cla_2/g0 cla_2/g1 0.26fF
C435 cla_0/nand_0/w_0_0# cla_0/n 0.04fF
C436 s4 sumffo_3/xor_0/inv_1/op 0.52fF
C437 sumffo_2/xor_0/inv_0/op sumffo_2/xor_0/w_n3_4# 0.06fF
C438 gnd ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C439 sumffo_3/xor_0/a_10_10# vdd 0.93fF
C440 cla_2/l cla_2/nor_0/w_0_0# 0.05fF
C441 nand_2/b sumffo_1/xor_0/inv_1/op 0.22fF
C442 cla_0/l nor_0/a 0.16fF
C443 ffipg_3/pggen_0/nor_0/a_13_6# ffipg_3/k 0.01fF
C444 cin sumffo_3/xor_0/a_10_10# 0.04fF
C445 ffipg_1/k vdd 0.36fF
C446 inv_2/in vdd 0.30fF
C447 inv_1/in nor_1/b 0.16fF
C448 cla_0/inv_0/in cla_0/g0 0.16fF
C449 inv_7/w_0_6# inv_7/op 0.03fF
C450 ffipg_1/k cin 0.06fF
C451 inv_2/in cin 0.13fF
C452 inv_8/w_0_6# vdd 0.15fF
C453 gnd inv_9/in 0.24fF
C454 cla_0/l cla_0/inv_0/in 0.14fF
C455 nand_2/b inv_2/w_0_6# 0.03fF
C456 gnd y2in 1.68fF
C457 cla_0/nor_0/w_0_0# vdd 0.31fF
C458 nand_2/b sumffo_2/c 0.06fF
C459 inv_8/w_0_6# cin 0.06fF
C460 x4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C461 y3in ffipg_2/pggen_0/xor_0/a_10_10# 0.12fF
C462 vdd nor_4/w_0_0# 0.15fF
C463 cla_0/nand_0/w_0_0# nand_2/b 0.05fF
C464 ffipg_3/pggen_0/xor_0/w_n3_4# ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C465 ffipg_1/k ffipg_1/pggen_0/xor_0/w_n3_4# 0.02fF
C466 inv_1/op sumffo_2/xor_0/inv_1/op 0.06fF
C467 cla_2/nand_0/w_0_0# cla_2/inv_0/op 0.06fF
C468 ffipg_0/pggen_0/xor_0/inv_0/op x1in 0.27fF
C469 x4in ffipg_3/pggen_0/xor_0/inv_1/op 0.06fF
C470 cla_2/g0 gnd 0.27fF
C471 cla_0/inv_0/in cla_0/inv_0/op 0.04fF
C472 inv_8/in vdd 0.30fF
C473 y3in ffipg_2/pggen_0/nand_0/w_0_0# 0.06fF
C474 ffipg_1/k y2in 0.07fF
C475 cla_2/g1 cla_2/inv_0/op 0.35fF
C476 gnd inv_5/in 0.19fF
C477 cin inv_8/in 0.13fF
C478 nor_3/b cla_2/n 0.41fF
C479 cla_2/p0 cla_1/inv_0/in 0.02fF
C480 sumffo_2/xor_0/inv_0/op vdd 0.15fF
C481 cla_1/nand_0/w_0_0# cla_1/n 0.04fF
C482 inv_7/w_0_6# vdd 0.15fF
C483 nor_2/b vdd 0.21fF
C484 ffipg_0/k sumffo_0/xor_0/w_n3_4# 0.06fF
C485 cin sumffo_2/xor_0/inv_0/op 0.06fF
C486 sumffo_0/xor_0/inv_1/op s1 0.52fF
C487 nor_4/w_0_0# inv_9/in 0.11fF
C488 vdd sumffo_2/xor_0/w_n3_4# 0.12fF
C489 cla_2/p0 ffipg_2/pggen_0/nand_0/w_0_0# 0.24fF
C490 gnd sumffo_0/xor_0/inv_0/op 0.21fF
C491 cin sumffo_2/xor_0/w_n3_4# 0.00fF
C492 vdd y1in 0.15fF
C493 gnd nor_3/b 0.10fF
C494 inv_7/op vdd 0.17fF
C495 inv_0/in nor_0/a 0.02fF
C496 sumffo_3/xor_0/inv_0/op vdd 0.15fF
C497 sumffo_0/xor_0/inv_1/op sumffo_0/xor_0/inv_1/w_0_6# 0.03fF
C498 ffipg_0/k sumffo_0/xor_0/inv_0/op 0.27fF
C499 sumffo_3/xor_0/w_n3_4# sumffo_3/xor_0/inv_1/op 0.06fF
C500 gnd inv_1/in 0.24fF
C501 ffipg_0/pggen_0/xor_0/inv_0/op ffipg_0/pggen_0/xor_0/inv_0/w_0_6# 0.03fF
C502 cin inv_7/op 0.31fF
C503 cla_2/p1 ffipg_3/pggen_0/nand_0/w_0_0# 0.24fF
C504 ffipg_3/k ffipg_3/pggen_0/xor_0/inv_1/op 0.52fF
C505 nor_3/w_0_0# inv_6/in 0.11fF
C506 gnd inv_0/op 0.10fF
C507 gnd sumffo_0/xor_0/inv_0/w_0_6# 0.02fF
C508 ffipg_0/k ffipg_0/pggen_0/xor_0/w_n3_4# 0.02fF
C509 ffipg_2/k x3in 0.46fF
C510 gnd cla_2/inv_0/op 0.10fF
C511 ffipg_0/k sumffo_0/xor_0/inv_0/w_0_6# 0.06fF
C512 nor_0/a x1in 0.22fF
C513 nand_2/b sumffo_1/xor_0/inv_0/op 0.20fF
C514 sumffo_1/xor_0/w_n3_4# vdd 0.12fF
C515 cla_0/n nor_1/b 0.36fF
C516 sumffo_1/xor_0/w_n3_4# cin 0.00fF
C517 gnd sumffo_3/xor_0/inv_1/op 0.20fF
C518 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/k 0.02fF
C519 ffipg_2/pggen_0/xor_0/inv_1/op vdd 0.15fF
C520 gnd cla_1/nand_0/w_0_0# 0.01fF
C521 cla_0/l inv_3/in 0.22fF
C522 y4in ffipg_3/pggen_0/nand_0/w_0_0# 0.06fF
C523 sumffo_3/xor_0/inv_0/w_0_6# sumffo_3/xor_0/inv_0/op 0.03fF
C524 cla_1/g0 vdd 0.55fF
C525 gnd x4in 0.31fF
C526 gnd cla_1/p0 0.68fF
C527 gnd y3in 1.68fF
C528 gnd sumffo_2/xor_0/inv_1/op 0.20fF
C529 cla_2/inv_0/in cla_2/nor_1/w_0_0# 0.05fF
C530 cla_1/nor_0/w_0_0# cla_1/l 0.05fF
C531 cin vdd 0.78fF
C532 y4in ffipg_3/pggen_0/xor_0/inv_1/op 0.22fF
C533 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# ffipg_1/pggen_0/xor_0/inv_0/op 0.03fF
C534 nand_2/b sumffo_1/xor_0/a_10_10# 0.12fF
C535 cla_0/l cla_2/l 0.37fF
C536 ffipg_3/k sumffo_3/xor_0/w_n3_4# 0.06fF
C537 sumffo_0/xor_0/a_10_10# s1 0.45fF
C538 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/k 0.06fF
C539 ffipg_2/pggen_0/xor_0/w_n3_4# x3in 0.06fF
C540 vdd inv_5/w_0_6# 0.15fF
C541 cla_2/g1 cla_2/p1 0.00fF
C542 cinbar inv_0/in 0.16fF
C543 cla_1/inv_0/in cla_1/inv_0/op 0.04fF
C544 gnd s3 0.14fF
C545 gnd cla_2/p0 0.68fF
C546 cla_0/n inv_3/w_0_6# 0.16fF
C547 ffipg_1/pggen_0/xor_0/w_n3_4# vdd 0.12fF
C548 nor_4/b inv_6/in 0.04fF
C549 ffipg_1/k cla_1/p0 0.05fF
C550 gnd cout 0.10fF
C551 cla_1/inv_0/in cla_1/nor_1/w_0_0# 0.05fF
C552 cla_1/g0 y2in 0.13fF
C553 sumffo_2/c ffipg_2/k 0.03fF
C554 ffipg_0/pggen_0/nand_0/w_0_0# y1in 0.06fF
C555 vdd inv_9/in 0.09fF
C556 ffipg_2/pggen_0/xor_0/inv_0/op x3in 0.27fF
C557 cla_1/p0 cla_0/nor_0/w_0_0# 0.06fF
C558 y2in vdd 0.15fF
C559 sumffo_3/xor_0/inv_0/w_0_6# vdd 0.09fF
C560 cla_0/l cla_0/inv_0/op 0.21fF
C561 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# y4in 0.23fF
C562 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# ffipg_0/pggen_0/xor_0/inv_1/op 0.03fF
C563 gnd ffipg_3/k 0.31fF
C564 x1in ffipg_0/pggen_0/xor_0/inv_1/op 0.06fF
C565 cla_2/g1 y4in 0.13fF
C566 nand_2/b inv_3/w_0_6# 0.06fF
C567 inv_1/op nor_1/w_0_0# 0.03fF
C568 gnd cla_0/n 0.61fF
C569 cla_2/g0 cla_1/g0 0.35fF
C570 y1in ffipg_0/pggen_0/xor_0/w_n3_4# 0.06fF
C571 gnd ffipg_0/pggen_0/xor_0/inv_0/op 0.17fF
C572 nand_2/b sumffo_1/xor_0/inv_1/w_0_6# 0.23fF
C573 gnd cla_2/p1 0.68fF
C574 ffipg_1/k ffipg_1/pggen_0/xor_0/a_10_10# 0.45fF
C575 sumffo_2/xor_0/a_10_10# sumffo_2/c 0.12fF
C576 ffipg_2/pggen_0/xor_0/inv_0/op ffipg_2/pggen_0/xor_0/w_n3_4# 0.06fF
C577 cla_2/g0 vdd 0.56fF
C578 ffipg_0/k ffipg_0/pggen_0/xor_0/inv_0/op 0.06fF
C579 y2in ffipg_1/pggen_0/xor_0/w_n3_4# 0.06fF
C580 ffipg_3/k sumffo_3/xor_0/a_10_10# 0.12fF
C581 ffipg_0/pggen_0/nor_0/w_0_0# x1in 0.06fF
C582 cla_1/inv_0/w_0_6# cla_1/inv_0/in 0.06fF
C583 inv_5/in vdd 0.30fF
C584 sumffo_2/xor_0/inv_0/w_0_6# inv_1/op 0.06fF
C585 cout nor_4/w_0_0# 0.03fF
C586 nor_3/w_0_0# cla_2/n 0.06fF
C587 cla_0/l inv_2/w_0_6# 0.06fF
C588 ffipg_3/pggen_0/xor_0/inv_0/op ffipg_3/pggen_0/xor_0/inv_1/op 0.08fF
C589 cla_0/l sumffo_2/c 0.04fF
C590 sumffo_2/xor_0/inv_1/w_0_6# vdd 0.06fF
C591 sumffo_0/xor_0/w_n3_4# vdd 0.12fF
C592 nor_1/w_0_0# nor_1/b 0.06fF
C593 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/inv_0/op 0.08fF
C594 cla_0/nand_0/w_0_0# cla_0/l 0.00fF
C595 ffipg_1/pggen_0/nor_0/w_0_0# x2in 0.06fF
C596 gnd nand_2/b 0.94fF
C597 sumffo_0/xor_0/w_n3_4# cin 0.06fF
C598 sumffo_3/xor_0/inv_0/op sumffo_3/xor_0/inv_1/op 0.08fF
C599 inv_5/in inv_5/w_0_6# 0.10fF
C600 ffipg_0/pggen_0/nand_0/w_0_0# vdd 0.10fF
C601 sumffo_2/xor_0/inv_1/op sumffo_2/xor_0/w_n3_4# 0.06fF
C602 sumffo_0/xor_0/inv_0/op vdd 0.15fF
C603 gnd y4in 1.66fF
C604 gnd cla_0/nand_0/a_13_n26# 0.00fF
C605 vdd ffipg_2/pggen_0/xor_0/inv_0/w_0_6# 0.09fF
C606 nor_3/b vdd 0.23fF
C607 sumffo_0/xor_0/inv_0/op cin 0.20fF
C608 inv_1/in vdd 0.09fF
C609 s3 sumffo_2/xor_0/inv_0/op 0.06fF
C610 cla_0/nand_0/w_0_0# cla_0/inv_0/op 0.06fF
C611 vdd ffipg_0/pggen_0/xor_0/w_n3_4# 0.12fF
C612 sumffo_1/xor_0/inv_0/w_0_6# sumffo_1/xor_0/inv_0/op 0.03fF
C613 gnd cla_1/inv_0/op 0.10fF
C614 inv_0/op vdd 0.17fF
C615 s3 sumffo_2/xor_0/w_n3_4# 0.02fF
C616 sumffo_0/xor_0/inv_0/w_0_6# vdd 0.09fF
C617 nor_3/b inv_5/w_0_6# 0.17fF
C618 inv_2/in nand_2/b 0.34fF
C619 nand_2/b ffipg_1/k 0.15fF
C620 cla_2/inv_0/op vdd 0.17fF
C621 ffipg_2/pggen_0/xor_0/a_10_10# ffipg_2/k 0.45fF
C622 gnd nor_0/a 0.23fF
C623 gnd cla_2/nand_0/a_13_n26# 0.01fF
C624 ffipg_0/k nor_0/a 0.05fF
C625 vdd sumffo_3/xor_0/inv_1/op 0.15fF
C626 ffipg_2/pggen_0/xor_0/inv_1/op y3in 0.22fF
C627 nor_4/a nor_4/b 0.42fF
C628 vdd ffipg_3/pggen_0/xor_0/w_n3_4# 0.12fF
C629 gnd cla_0/inv_0/in 0.30fF
C630 cla_1/nand_0/w_0_0# vdd 0.10fF
C631 cla_1/g0 cla_1/p0 0.07fF
C632 cla_1/g0 cla_0/nor_1/w_0_0# 0.02fF
C633 cin sumffo_3/xor_0/inv_1/op 0.04fF
C634 x4in vdd 0.93fF
C635 cla_1/p0 vdd 0.43fF
C636 ffipg_3/k sumffo_3/xor_0/inv_0/op 0.20fF
C637 cla_0/nor_1/w_0_0# vdd 0.31fF
C638 y3in vdd 0.15fF
C639 ffipg_2/pggen_0/xor_0/inv_1/op ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.03fF
C640 sumffo_2/xor_0/inv_1/op vdd 0.15fF
C641 vdd ffipg_2/pggen_0/nor_0/w_0_0# 0.11fF
C642 ffipg_0/pggen_0/xor_0/inv_0/op y1in 0.20fF
C643 ffipg_1/k nor_0/a 0.06fF
C644 cin sumffo_2/xor_0/inv_1/op 0.04fF
C645 gnd nor_4/b 0.10fF
C646 gnd ffipg_3/pggen_0/xor_0/inv_0/op 0.21fF
C647 vdd ffipg_2/pggen_0/xor_0/inv_1/w_0_6# 0.06fF
C648 cla_2/g1 cla_2/inv_0/in 0.04fF
C649 cla_2/p0 cla_1/g0 0.36fF
C650 ffipg_2/pggen_0/nor_0/a_13_6# ffipg_2/k 0.01fF
C651 ffipg_1/k ffipg_1/pggen_0/nor_0/a_13_6# 0.01fF
C652 cla_2/p0 vdd 0.43fF
C653 cla_0/nor_0/w_0_0# nor_0/a 0.06fF
C654 ffipg_2/pggen_0/xor_0/w_n3_4# ffipg_2/pggen_0/xor_0/a_10_10# 0.16fF
C655 nor_3/b inv_5/in 0.04fF
C656 sumffo_0/xor_0/inv_0/op sumffo_0/xor_0/w_n3_4# 0.06fF
C657 inv_3/w_0_6# cla_1/l 0.06fF
C658 ffipg_3/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C659 ffipg_3/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C660 ffipg_3/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C661 ffipg_3/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C662 ffipg_3/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C663 ffipg_3/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C664 ffipg_3/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C665 y4in Gnd 2.72fF
C666 x4in Gnd 2.80fF
C667 ffipg_3/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C668 ffipg_2/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C669 ffipg_2/k Gnd 1.51fF
C670 ffipg_2/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C671 ffipg_2/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C672 ffipg_2/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C673 ffipg_2/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C674 ffipg_2/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C675 ffipg_2/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C676 y3in Gnd 2.72fF
C677 x3in Gnd 2.80fF
C678 ffipg_2/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C679 ffipg_1/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C680 ffipg_1/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C681 ffipg_1/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C682 ffipg_1/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C683 ffipg_1/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C684 ffipg_1/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C685 ffipg_1/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C686 y2in Gnd 2.72fF
C687 x2in Gnd 2.80fF
C688 ffipg_1/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C689 cout Gnd 0.19fF
C690 inv_9/in Gnd 0.23fF
C691 nor_4/w_0_0# Gnd 1.81fF
C692 ffipg_0/pggen_0/nor_0/w_0_0# Gnd 1.23fF
C693 ffipg_0/pggen_0/xor_0/a_10_10# Gnd 0.01fF
C694 ffipg_0/pggen_0/xor_0/w_n3_4# Gnd 1.14fF
C695 ffipg_0/pggen_0/xor_0/inv_1/op Gnd 0.49fF
C696 ffipg_0/pggen_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C697 ffipg_0/pggen_0/xor_0/inv_0/op Gnd 0.50fF
C698 ffipg_0/pggen_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C699 y1in Gnd 2.72fF
C700 x1in Gnd 2.80fF
C701 ffipg_0/pggen_0/nand_0/w_0_0# Gnd 0.82fF
C702 nor_4/a Gnd 0.59fF
C703 inv_8/in Gnd 0.22fF
C704 inv_8/w_0_6# Gnd 1.40fF
C705 inv_7/in Gnd 0.22fF
C706 inv_7/w_0_6# Gnd 1.40fF
C707 nor_4/b Gnd 0.32fF
C708 nor_3/b Gnd 0.77fF
C709 inv_5/in Gnd 0.22fF
C710 inv_5/w_0_6# Gnd 1.40fF
C711 cla_2/n Gnd 0.36fF
C712 inv_6/in Gnd 0.23fF
C713 nor_3/w_0_0# Gnd 1.81fF
C714 vdd Gnd 8.88fF
C715 cla_1/n Gnd 0.36fF
C716 inv_4/in Gnd 0.23fF
C717 nor_2/w_0_0# Gnd 1.81fF
C718 cla_0/n Gnd 1.34fF
C719 nor_2/b Gnd 0.82fF
C720 inv_3/in Gnd 0.22fF
C721 inv_3/w_0_6# Gnd 1.40fF
C722 cinbar Gnd 1.21fF
C723 nor_0/a Gnd 2.07fF
C724 nor_1/b Gnd 1.05fF
C725 inv_2/in Gnd 0.22fF
C726 inv_2/w_0_6# Gnd 1.40fF
C727 inv_1/in Gnd 0.23fF
C728 nor_1/w_0_0# Gnd 1.81fF
C729 inv_0/in Gnd 0.23fF
C730 s4 Gnd 0.07fF
C731 sumffo_3/xor_0/a_10_10# Gnd 0.01fF
C732 sumffo_3/xor_0/w_n3_4# Gnd 1.14fF
C733 sumffo_3/xor_0/inv_1/op Gnd 0.49fF
C734 ffipg_3/k Gnd 2.89fF
C735 sumffo_3/xor_0/inv_1/w_0_6# Gnd 0.58fF
C736 sumffo_3/xor_0/inv_0/op Gnd 0.50fF
C737 inv_4/op Gnd 1.37fF
C738 sumffo_3/xor_0/inv_0/w_0_6# Gnd 0.58fF
C739 s2 Gnd 0.07fF
C740 sumffo_1/xor_0/a_10_10# Gnd 0.01fF
C741 sumffo_1/xor_0/w_n3_4# Gnd 1.14fF
C742 sumffo_1/xor_0/inv_1/op Gnd 0.49fF
C743 nand_2/b Gnd 2.36fF
C744 sumffo_1/xor_0/inv_1/w_0_6# Gnd 0.58fF
C745 sumffo_1/xor_0/inv_0/op Gnd 0.50fF
C746 ffipg_1/k Gnd 2.78fF
C747 sumffo_1/xor_0/inv_0/w_0_6# Gnd 0.58fF
C748 s3 Gnd 0.07fF
C749 sumffo_2/xor_0/a_10_10# Gnd 0.01fF
C750 sumffo_2/xor_0/w_n3_4# Gnd 1.14fF
C751 sumffo_2/xor_0/inv_1/op Gnd 0.49fF
C752 sumffo_2/c Gnd 1.92fF
C753 sumffo_2/xor_0/inv_1/w_0_6# Gnd 0.58fF
C754 sumffo_2/xor_0/inv_0/op Gnd 0.50fF
C755 inv_1/op Gnd 1.30fF
C756 sumffo_2/xor_0/inv_0/w_0_6# Gnd 0.58fF
C757 s1 Gnd 0.07fF
C758 sumffo_0/xor_0/a_10_10# Gnd 0.01fF
C759 sumffo_0/xor_0/w_n3_4# Gnd 1.14fF
C760 gnd Gnd 23.13fF
C761 sumffo_0/xor_0/inv_1/op Gnd 0.49fF
C762 cin Gnd 7.80fF
C763 sumffo_0/xor_0/inv_1/w_0_6# Gnd 0.58fF
C764 sumffo_0/xor_0/inv_0/op Gnd 0.50fF
C765 ffipg_0/k Gnd 1.49fF
C766 sumffo_0/xor_0/inv_0/w_0_6# Gnd 0.58fF
C767 cla_2/p1 Gnd 1.09fF
C768 cla_2/nor_1/w_0_0# Gnd 1.23fF
C769 cla_2/nor_0/w_0_0# Gnd 1.23fF
C770 cla_2/inv_0/in Gnd 0.27fF
C771 cla_2/inv_0/w_0_6# Gnd 0.58fF
C772 cla_2/g1 Gnd 0.59fF
C773 cla_2/inv_0/op Gnd 0.26fF
C774 cla_2/nand_0/w_0_0# Gnd 0.82fF
C775 cla_2/p0 Gnd 0.38fF
C776 cla_1/nor_1/w_0_0# Gnd 1.23fF
C777 cla_1/l Gnd 0.30fF
C778 cla_1/nor_0/w_0_0# Gnd 1.23fF
C779 cla_1/inv_0/in Gnd 0.27fF
C780 cla_1/inv_0/w_0_6# Gnd 0.58fF
C781 cla_2/g0 Gnd 1.58fF
C782 cla_1/inv_0/op Gnd 0.26fF
C783 cla_1/nand_0/w_0_0# Gnd 0.82fF
C784 inv_7/op Gnd 0.26fF
C785 cla_1/p0 Gnd 2.28fF
C786 cla_0/nor_1/w_0_0# Gnd 1.23fF
C787 cla_0/l Gnd 0.45fF
C788 cla_0/nor_0/w_0_0# Gnd 1.23fF
C789 cla_0/inv_0/in Gnd 0.27fF
C790 cla_0/inv_0/w_0_6# Gnd 0.58fF
C791 cla_1/g0 Gnd 1.49fF
C792 cla_0/inv_0/op Gnd 0.26fF
C793 cla_0/nand_0/w_0_0# Gnd 0.82fF
C794 cla_2/l Gnd 0.25fF
C795 cla_0/g0 Gnd 1.40fF
C796 inv_0/op Gnd 0.23fF
C797 nor_0/w_0_0# Gnd 2.63fF
